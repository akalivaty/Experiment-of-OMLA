//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  OAI211_X1 g007(.A(KEYINPUT23), .B(new_n204), .C1(new_n206), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n209), .A2(new_n213), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(KEYINPUT25), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n235));
  OAI211_X1 g034(.A(KEYINPUT28), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT28), .A4(new_n233), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n207), .A2(new_n204), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(KEYINPUT26), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(KEYINPUT26), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n210), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n214), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  INV_X1    g050(.A(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G113gat), .ZN(new_n255));
  INV_X1    g054(.A(G113gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT1), .B(G127gat), .C1(new_n255), .C2(new_n257), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n252), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G120gat), .ZN(new_n263));
  OAI21_X1  g062(.A(G127gat), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n258), .A2(new_n259), .A3(new_n253), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n250), .A2(new_n251), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n251), .B1(new_n250), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n250), .A2(new_n267), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n203), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT32), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT34), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n244), .A2(new_n214), .A3(new_n248), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n225), .A2(new_n226), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n221), .B1(new_n278), .B2(new_n223), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n279), .A2(new_n230), .B1(new_n220), .B2(new_n221), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n267), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT67), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n250), .A2(new_n251), .A3(new_n267), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n271), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n203), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n284), .A2(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n287), .B1(new_n286), .B2(KEYINPUT32), .ZN(new_n292));
  AOI211_X1 g091(.A(new_n273), .B(KEYINPUT34), .C1(new_n284), .C2(new_n285), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT68), .B(G71gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n272), .B2(KEYINPUT33), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n291), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n291), .B2(new_n294), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n202), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n292), .A2(new_n293), .A3(new_n289), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n290), .B1(new_n274), .B2(new_n288), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n294), .A3(new_n300), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(KEYINPUT36), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  NOR2_X1   g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316));
  NAND2_X1  g115(.A1(G211gat), .A2(G218gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(KEYINPUT69), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n275), .B2(new_n280), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n232), .B2(new_n249), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n322), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n325), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(new_n250), .B2(new_n323), .ZN(new_n331));
  INV_X1    g130(.A(new_n322), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n331), .A2(new_n332), .A3(new_n327), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n309), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G8gat), .B(G36gat), .Z(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(G64gat), .ZN(new_n336));
  INV_X1    g135(.A(G92gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT72), .Z(new_n339));
  NAND3_X1  g138(.A1(new_n326), .A2(new_n322), .A3(new_n328), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n332), .B1(new_n331), .B2(new_n327), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT71), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n334), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n338), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n352));
  OAI21_X1  g151(.A(G148gat), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G141gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(G148gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n360), .B2(KEYINPUT2), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT2), .ZN(new_n362));
  INV_X1    g161(.A(G148gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G141gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n355), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n358), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(new_n359), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n357), .A2(new_n361), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n262), .A2(new_n266), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n262), .A2(new_n368), .A3(KEYINPUT75), .A4(new_n266), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT74), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n368), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n368), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n267), .A3(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n369), .A2(new_n374), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n375), .A2(new_n378), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n368), .B1(new_n262), .B2(new_n266), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(new_n377), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n371), .B2(new_n372), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n391), .A2(KEYINPUT76), .A3(new_n378), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT5), .B(new_n385), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n374), .B1(new_n371), .B2(new_n372), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT78), .B1(new_n369), .B2(KEYINPUT4), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI211_X1 g201(.A(KEYINPUT78), .B(new_n374), .C1(new_n371), .C2(new_n372), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n404), .A3(new_n378), .ZN(new_n405));
  OR3_X1    g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n393), .A2(new_n399), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n399), .B1(new_n393), .B2(new_n406), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n389), .A2(new_n386), .A3(new_n377), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT76), .B1(new_n391), .B2(new_n378), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n404), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(new_n385), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n417), .A2(new_n399), .A3(new_n409), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n350), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT31), .B(G50gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G106gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G22gat), .B(G78gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT80), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n322), .B1(new_n323), .B2(new_n382), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n311), .A2(new_n318), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n311), .A2(new_n318), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n323), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n368), .B1(new_n431), .B2(new_n381), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n427), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n319), .B2(new_n321), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n379), .B1(new_n434), .B2(KEYINPUT3), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n382), .A2(new_n323), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n332), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n425), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n424), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n439), .A3(new_n424), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n422), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n442), .ZN(new_n444));
  INV_X1    g243(.A(new_n422), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n444), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n420), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n422), .A3(new_n442), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n445), .B1(new_n444), .B2(new_n440), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT81), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n303), .A2(new_n308), .B1(new_n419), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n389), .A2(new_n377), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n400), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(new_n383), .C1(new_n400), .C2(new_n401), .ZN(new_n459));
  AOI211_X1 g258(.A(new_n455), .B(new_n456), .C1(new_n459), .C2(new_n377), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n455), .A3(new_n377), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n399), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n454), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT40), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n417), .B2(new_n399), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n411), .A2(KEYINPUT83), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n454), .B(new_n469), .C1(new_n460), .C2(new_n462), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n464), .A2(new_n468), .A3(new_n349), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n408), .B1(new_n417), .B2(new_n399), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n393), .A2(new_n406), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT83), .B1(new_n473), .B2(new_n398), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n465), .B(new_n399), .C1(new_n393), .C2(new_n406), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n411), .A2(new_n408), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT84), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(KEYINPUT37), .C1(KEYINPUT84), .C2(new_n341), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  OR3_X1    g279(.A1(new_n329), .A2(new_n333), .A3(KEYINPUT37), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n339), .A4(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n482), .A2(new_n345), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n476), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n334), .A2(KEYINPUT37), .A3(new_n342), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n338), .A3(new_n481), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT38), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n486), .B2(KEYINPUT38), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n453), .B(new_n471), .C1(new_n484), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n443), .A2(new_n446), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n301), .A2(new_n302), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n349), .B1(new_n476), .B2(new_n477), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT35), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n306), .A2(new_n453), .A3(new_n307), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT35), .B1(new_n497), .B2(new_n419), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n452), .A2(new_n491), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500));
  INV_X1    g299(.A(G211gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G57gat), .B(G64gat), .Z(new_n504));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505));
  INV_X1    g304(.A(G71gat), .ZN(new_n506));
  INV_X1    g305(.A(G78gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n509), .A2(new_n510), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n510), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n516), .A3(new_n508), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT88), .B1(new_n517), .B2(new_n511), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT21), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n253), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n515), .A2(new_n518), .ZN(new_n522));
  OAI21_X1  g321(.A(G127gat), .B1(new_n522), .B2(KEYINPUT21), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G1gat), .B2(new_n525), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n519), .B2(new_n520), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n534));
  XNOR2_X1  g333(.A(G155gat), .B(G183gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n534), .B(new_n535), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n523), .A3(new_n521), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n533), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n533), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n503), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n538), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n531), .B1(new_n523), .B2(new_n521), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n533), .A2(new_n537), .A3(new_n538), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n502), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G162gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n551), .B2(KEYINPUT7), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT7), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n560), .B2(new_n337), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G99gat), .B(G106gat), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n565), .A3(new_n561), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G43gat), .B(G50gat), .Z(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  INV_X1    g368(.A(G36gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT14), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n572), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n574), .A2(G29gat), .A3(G36gat), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(new_n572), .B2(new_n571), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n568), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n568), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT17), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n568), .ZN(new_n585));
  INV_X1    g384(.A(new_n580), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n582), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n567), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n581), .A2(new_n583), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n564), .A3(new_n566), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G134gat), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n591), .A2(new_n594), .A3(new_n252), .A4(new_n592), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n596), .B2(new_n597), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n550), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n549), .A3(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n499), .A2(new_n547), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT87), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n584), .A2(new_n590), .A3(new_n530), .ZN(new_n609));
  INV_X1    g408(.A(new_n530), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n593), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT86), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n608), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT18), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n530), .B1(new_n581), .B2(new_n583), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n612), .B(KEYINPUT13), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT18), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n613), .B2(new_n608), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n616), .B(new_n620), .C1(new_n615), .C2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G197gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT11), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n207), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n615), .A2(new_n622), .ZN(new_n630));
  INV_X1    g429(.A(new_n628), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n620), .A4(new_n616), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n566), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n565), .B1(new_n558), .B2(new_n561), .ZN(new_n637));
  OAI22_X1  g436(.A1(new_n636), .A2(new_n637), .B1(new_n515), .B2(new_n518), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n562), .A2(KEYINPUT91), .A3(new_n563), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n512), .A2(new_n514), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n558), .A2(new_n561), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n522), .A2(KEYINPUT10), .A3(new_n564), .A4(new_n566), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n645), .A2(KEYINPUT92), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT92), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n635), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n635), .B1(new_n638), .B2(new_n643), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n204), .ZN(new_n653));
  INV_X1    g452(.A(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n649), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n645), .A2(new_n646), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n635), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n651), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n655), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n634), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n607), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n412), .A2(new_n418), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT93), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT94), .B(G1gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  NAND3_X1  g468(.A1(new_n607), .A2(new_n663), .A3(new_n349), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n607), .A2(KEYINPUT95), .A3(new_n663), .A4(new_n349), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n672), .B(KEYINPUT96), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT97), .B1(new_n677), .B2(G8gat), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n681), .B(new_n529), .C1(new_n675), .C2(new_n676), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n673), .B(new_n679), .C1(new_n680), .C2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(G15gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n303), .A2(new_n308), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n664), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n664), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n301), .A2(new_n302), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n684), .B2(new_n689), .ZN(G1326gat));
  INV_X1    g489(.A(new_n451), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n664), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n606), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n499), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n491), .A2(new_n452), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n496), .A2(new_n498), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n606), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n634), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n547), .B(KEYINPUT98), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n662), .B(KEYINPUT99), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT100), .B1(new_n706), .B2(new_n666), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n708));
  INV_X1    g507(.A(new_n666), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n702), .A2(new_n708), .A3(new_n709), .A4(new_n705), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(G29gat), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n699), .A2(new_n606), .ZN(new_n712));
  INV_X1    g511(.A(new_n547), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n714), .A2(new_n569), .A3(new_n709), .A4(new_n663), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(G1328gat));
  NAND4_X1  g516(.A1(new_n714), .A2(new_n570), .A3(new_n663), .A4(new_n349), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n718), .A2(new_n721), .A3(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n718), .B2(KEYINPUT46), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n706), .B2(new_n350), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n663), .ZN(new_n728));
  INV_X1    g527(.A(new_n688), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n685), .A2(new_n727), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n702), .A2(new_n705), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1330gat));
  NOR3_X1   g535(.A1(new_n728), .A2(G50gat), .A3(new_n691), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G50gat), .B1(new_n706), .B2(new_n453), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT48), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n702), .A2(new_n451), .A3(new_n705), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n737), .B1(G50gat), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g542(.A1(new_n633), .A2(new_n547), .A3(new_n606), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n704), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT104), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n699), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n709), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g549(.A(new_n350), .B(new_n747), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1333gat));
  NOR3_X1   g552(.A1(new_n747), .A2(new_n506), .A3(new_n685), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n688), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n506), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g556(.A1(new_n747), .A2(new_n691), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT105), .B(G78gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1335gat));
  AOI21_X1  g559(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n713), .A2(new_n633), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n766), .A2(new_n560), .A3(new_n709), .A4(new_n662), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n696), .A2(new_n701), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n762), .A2(new_n662), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g572(.A(KEYINPUT106), .B(new_n770), .C1(new_n696), .C2(new_n701), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n666), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n776), .B2(new_n560), .ZN(G1336gat));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n769), .A2(new_n771), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n778), .B(G92gat), .C1(new_n779), .C2(new_n350), .ZN(new_n780));
  INV_X1    g579(.A(new_n704), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n350), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n337), .B(new_n782), .C1(new_n783), .C2(new_n763), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n780), .B(new_n784), .C1(new_n785), .C2(new_n778), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n349), .B1(new_n772), .B2(new_n774), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(G92gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n778), .ZN(G1337gat));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n688), .A2(new_n791), .A3(new_n662), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT108), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n766), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n685), .B1(new_n773), .B2(new_n775), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n791), .ZN(G1338gat));
  INV_X1    g595(.A(G106gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n453), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n766), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G106gat), .B1(new_n779), .B2(new_n453), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n798), .ZN(new_n803));
  AOI211_X1 g602(.A(G106gat), .B(new_n803), .C1(new_n764), .C2(new_n765), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n451), .B1(new_n772), .B2(new_n774), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n802), .B1(new_n806), .B2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(new_n662), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n634), .A2(new_n695), .A3(new_n809), .A4(new_n713), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n744), .A2(new_n812), .A3(new_n809), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n815));
  INV_X1    g614(.A(new_n635), .ZN(new_n816));
  AOI211_X1 g615(.A(KEYINPUT54), .B(new_n816), .C1(new_n645), .C2(new_n646), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n817), .B2(new_n656), .ZN(new_n818));
  OAI211_X1 g617(.A(KEYINPUT111), .B(new_n655), .C1(new_n659), .C2(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n645), .A2(new_n816), .A3(new_n646), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n649), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n633), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n657), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n612), .B1(new_n609), .B2(new_n611), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n611), .A2(new_n617), .A3(new_n619), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(KEYINPUT113), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n830), .B2(new_n829), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n831), .A2(KEYINPUT113), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n627), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n632), .A2(new_n835), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n826), .A2(new_n828), .B1(new_n809), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n632), .A2(KEYINPUT114), .A3(new_n835), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT114), .B1(new_n632), .B2(new_n835), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT55), .B1(new_n820), .B2(new_n822), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n828), .A2(new_n695), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n837), .A2(new_n695), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n814), .B1(new_n843), .B2(new_n703), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n666), .A2(new_n349), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n493), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n256), .A3(new_n633), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n729), .A2(new_n451), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n634), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(G1340gat));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n254), .A3(new_n662), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n850), .B2(new_n781), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n847), .B2(new_n713), .ZN(new_n856));
  INV_X1    g655(.A(new_n703), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n850), .A2(new_n253), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n847), .A2(new_n252), .A3(new_n606), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n850), .B2(new_n695), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n863), .A3(new_n252), .A4(new_n606), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n811), .A2(new_n813), .ZN(new_n866));
  INV_X1    g665(.A(new_n838), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n839), .A2(new_n840), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n842), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n828), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n823), .A2(new_n824), .B1(new_n629), .B2(new_n632), .ZN(new_n871));
  INV_X1    g670(.A(new_n836), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n870), .A2(new_n871), .B1(new_n662), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(new_n606), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n866), .B1(new_n874), .B2(new_n547), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n691), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n844), .A2(new_n877), .A3(new_n492), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n845), .A2(new_n685), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n876), .A2(new_n878), .A3(new_n633), .A4(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n837), .A2(new_n695), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n713), .B1(new_n884), .B2(new_n869), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n451), .B1(new_n885), .B2(new_n866), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n886), .B2(KEYINPUT57), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(KEYINPUT116), .A3(new_n633), .A4(new_n878), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n351), .A2(new_n352), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n844), .A2(new_n492), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n354), .A3(new_n633), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n894), .A2(new_n897), .A3(new_n354), .A4(new_n633), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n874), .A2(new_n857), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n453), .B1(new_n899), .B2(new_n814), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n354), .A3(new_n880), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT115), .B1(new_n901), .B2(new_n634), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n881), .A2(new_n890), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT58), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n896), .A2(new_n905), .ZN(G1344gat));
  NAND3_X1  g705(.A1(new_n894), .A2(new_n363), .A3(new_n662), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n878), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n809), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(KEYINPUT59), .A3(new_n363), .ZN(new_n910));
  XOR2_X1   g709(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n911));
  NAND2_X1  g710(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n810), .B(KEYINPUT118), .Z(new_n913));
  OAI211_X1 g712(.A(new_n877), .B(new_n451), .C1(new_n913), .C2(new_n885), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n912), .A2(new_n662), .A3(new_n914), .A4(new_n880), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n910), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(G155gat), .B1(new_n894), .B2(new_n713), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n887), .A2(new_n878), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n703), .A2(G155gat), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT119), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n908), .B2(new_n695), .ZN(new_n923));
  INV_X1    g722(.A(G162gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n894), .A2(new_n924), .A3(new_n606), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(KEYINPUT120), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(KEYINPUT120), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1347gat));
  NAND4_X1  g727(.A1(new_n844), .A2(new_n666), .A3(new_n349), .A4(new_n849), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n634), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n709), .B1(new_n899), .B2(new_n814), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n493), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n349), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n633), .B1(new_n206), .B2(new_n208), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  NOR3_X1   g734(.A1(new_n929), .A2(new_n204), .A3(new_n781), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n662), .A3(new_n349), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n204), .ZN(G1349gat));
  NAND4_X1  g737(.A1(new_n932), .A2(new_n238), .A3(new_n349), .A4(new_n713), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n929), .B2(new_n857), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT121), .B(KEYINPUT60), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OR2_X1    g740(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n942));
  NAND2_X1  g741(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n943));
  AND4_X1   g742(.A1(new_n942), .A2(new_n939), .A3(new_n943), .A4(new_n940), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n941), .A2(new_n944), .ZN(G1350gat));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n947));
  OAI211_X1 g746(.A(G190gat), .B(new_n947), .C1(new_n929), .C2(new_n695), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n233), .A3(new_n349), .A4(new_n606), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n349), .A3(new_n606), .A4(new_n849), .ZN(new_n952));
  INV_X1    g751(.A(new_n949), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n952), .A2(G190gat), .A3(new_n947), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n950), .A2(new_n957), .A3(new_n951), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1351gat));
  AND2_X1   g758(.A1(new_n912), .A2(new_n914), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n666), .A2(new_n349), .A3(new_n685), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT124), .Z(new_n963));
  NAND4_X1  g762(.A1(new_n960), .A2(new_n961), .A3(new_n633), .A4(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n963), .A2(new_n912), .A3(new_n633), .A4(new_n914), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(G197gat), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n900), .A2(new_n962), .ZN(new_n968));
  INV_X1    g767(.A(G197gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n633), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n970), .ZN(G1352gat));
  NAND2_X1  g770(.A1(new_n960), .A2(new_n963), .ZN(new_n972));
  OAI21_X1  g771(.A(G204gat), .B1(new_n972), .B2(new_n781), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n968), .A2(new_n654), .A3(new_n662), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n977), .B1(KEYINPUT126), .B2(new_n975), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n974), .A2(new_n979), .A3(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n973), .A2(new_n978), .A3(new_n980), .ZN(G1353gat));
  NAND2_X1  g780(.A1(new_n912), .A2(new_n914), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n962), .A2(new_n713), .ZN(new_n983));
  OAI21_X1  g782(.A(G211gat), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n984), .A2(KEYINPUT63), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(KEYINPUT63), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n501), .A3(new_n713), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n968), .A2(KEYINPUT127), .A3(new_n501), .A4(new_n713), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n985), .A2(new_n986), .A3(new_n991), .ZN(G1354gat));
  INV_X1    g791(.A(G218gat), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n972), .A2(new_n993), .A3(new_n695), .ZN(new_n994));
  AOI21_X1  g793(.A(G218gat), .B1(new_n968), .B2(new_n606), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


