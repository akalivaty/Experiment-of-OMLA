//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(new_n206), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NOR3_X1   g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n210), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n212), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n213), .B2(new_n218), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G77), .A2(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G116), .ZN(new_n224));
  INV_X1    g0024(.A(G270), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G97), .A2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G87), .A2(G250), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n230), .B1(new_n201), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(G107), .B2(G264), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(new_n216), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n221), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n231), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  INV_X1    g0040(.A(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n225), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n224), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  OAI21_X1  g0055(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR3_X1   g0059(.A1(KEYINPUT69), .A2(G20), .A3(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n210), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n267), .B2(KEYINPUT8), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n256), .B1(new_n257), .B2(new_n261), .C1(new_n262), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n211), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  INV_X1    g0072(.A(G13), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n273), .A2(new_n210), .A3(G1), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n269), .A2(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n271), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n214), .A2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G223), .A3(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G222), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n291), .B1(new_n253), .B2(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n285), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n283), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n241), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n282), .A2(KEYINPUT9), .B1(new_n300), .B2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n275), .A2(new_n281), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n301), .A2(new_n309), .A3(new_n303), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n300), .A2(G179), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n300), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n304), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n274), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G77), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G20), .A2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT15), .B(G87), .Z(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n319), .B1(new_n261), .B2(new_n320), .C1(new_n322), .C2(new_n262), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n323), .B2(new_n271), .ZN(new_n324));
  INV_X1    g0124(.A(new_n271), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G77), .A3(new_n278), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n326), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n318), .B(new_n330), .C1(new_n323), .C2(new_n271), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n290), .A2(G238), .A3(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n290), .A2(G232), .A3(new_n292), .ZN(new_n335));
  INV_X1    g0135(.A(G107), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n290), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n296), .ZN(new_n338));
  INV_X1    g0138(.A(new_n285), .ZN(new_n339));
  INV_X1    g0139(.A(new_n299), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G244), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n313), .ZN(new_n343));
  INV_X1    g0143(.A(new_n342), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n333), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n316), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  OAI211_X1 g0151(.A(G226), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(G223), .B(new_n292), .C1(new_n350), .C2(new_n351), .ZN(new_n353));
  INV_X1    g0153(.A(G87), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n352), .B(new_n353), .C1(new_n287), .C2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n285), .B1(new_n355), .B2(new_n296), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n340), .A2(G232), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G190), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n360), .B1(new_n356), .B2(new_n357), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n359), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n288), .A2(new_n210), .A3(new_n289), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n350), .A2(new_n351), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n205), .B(new_n203), .C1(new_n267), .C2(new_n202), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(G68), .B1(new_n374), .B2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(new_n261), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G159), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n367), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n371), .B2(new_n210), .ZN(new_n379));
  NOR4_X1   g0179(.A1(new_n350), .A2(new_n351), .A3(new_n369), .A4(G20), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n374), .A2(G20), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n367), .A4(new_n377), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n271), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n268), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n280), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n268), .A2(new_n274), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT17), .B1(new_n366), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n358), .A2(KEYINPUT76), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n365), .A3(new_n361), .ZN(new_n392));
  INV_X1    g0192(.A(new_n359), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n381), .A2(new_n377), .A3(new_n382), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n383), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n271), .B1(new_n386), .B2(new_n280), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n394), .A2(new_n398), .A3(new_n399), .A4(new_n388), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n390), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n362), .A2(new_n363), .A3(G169), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n398), .B2(new_n388), .ZN(new_n403));
  INV_X1    g0203(.A(new_n358), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n345), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT18), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n364), .A2(new_n313), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n389), .A2(new_n407), .A3(KEYINPUT18), .A4(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n401), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n331), .A2(KEYINPUT71), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT72), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n342), .A2(G200), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n329), .A2(new_n332), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT73), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n344), .A2(G190), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT73), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n416), .A2(new_n419), .A3(new_n423), .A4(new_n417), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G97), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n426), .B1(new_n287), .B2(new_n427), .C1(new_n293), .C2(new_n241), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n285), .B1(new_n428), .B2(new_n296), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n340), .A2(G238), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g0235(.A(new_n432), .ZN(new_n436));
  INV_X1    g0236(.A(new_n433), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(G179), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(G169), .C1(new_n432), .C2(new_n433), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n214), .A2(new_n202), .A3(G13), .A4(G20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n443));
  XOR2_X1   g0243(.A(new_n443), .B(KEYINPUT12), .Z(new_n444));
  NAND3_X1  g0244(.A1(new_n325), .A2(G68), .A3(new_n278), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g0246(.A(new_n446), .B(KEYINPUT75), .Z(new_n447));
  NOR2_X1   g0247(.A1(new_n261), .A2(new_n272), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n262), .A2(new_n253), .B1(new_n210), .B2(G68), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n271), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT11), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n436), .A2(G190), .A3(new_n437), .ZN(new_n455));
  OAI21_X1  g0255(.A(G200), .B1(new_n432), .B2(new_n433), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n425), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n349), .A2(new_n412), .A3(new_n413), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n276), .B1(G1), .B2(new_n287), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n336), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n274), .A2(new_n336), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT25), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n210), .B(G87), .C1(new_n350), .C2(new_n351), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT22), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n290), .A2(new_n468), .A3(new_n210), .A4(G87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n210), .A2(G107), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT23), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n473));
  XOR2_X1   g0273(.A(new_n473), .B(KEYINPUT84), .Z(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n470), .A2(new_n477), .A3(new_n474), .A4(new_n472), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n463), .B(new_n465), .C1(new_n479), .C2(new_n271), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n481));
  OAI211_X1 g0281(.A(G250), .B(new_n292), .C1(new_n350), .C2(new_n351), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G294), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n296), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT85), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G41), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n214), .B(G45), .C1(new_n488), .C2(KEYINPUT5), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT79), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G1), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G41), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT79), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n488), .A2(KEYINPUT5), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(G274), .A3(new_n298), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n296), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n488), .A2(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n214), .A2(G45), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n490), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n495), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G264), .A3(new_n298), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n487), .A2(new_n499), .A3(new_n500), .A4(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G190), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n485), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n506), .A2(new_n485), .A3(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(G200), .B1(new_n513), .B2(new_n499), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n480), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n505), .A2(G257), .A3(new_n298), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n499), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(new_n292), .C1(new_n350), .C2(new_n351), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n296), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n499), .A2(KEYINPUT80), .A3(new_n516), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n519), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n528), .A2(new_n516), .A3(new_n499), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G190), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n373), .A2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n336), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n427), .A2(new_n336), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n534), .B(new_n540), .C1(new_n253), .C2(new_n261), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n271), .B1(new_n427), .B2(new_n274), .ZN(new_n542));
  INV_X1    g0342(.A(new_n462), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G97), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n531), .A2(new_n533), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n544), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n528), .A2(new_n516), .A3(new_n499), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n313), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n519), .A2(new_n345), .A3(new_n528), .A4(new_n529), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n515), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n274), .A2(new_n224), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n543), .A2(G116), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n526), .B(new_n210), .C1(G33), .C2(new_n427), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(new_n271), .C1(new_n210), .C2(G116), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT83), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n552), .B(new_n553), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(new_n292), .C1(new_n350), .C2(new_n351), .ZN(new_n561));
  OAI211_X1 g0361(.A(G264), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n562));
  INV_X1    g0362(.A(G303), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n290), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n296), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n505), .A2(G270), .A3(new_n298), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n499), .A2(G179), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n560), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n499), .A2(new_n565), .A3(new_n566), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n572), .C1(new_n302), .C2(new_n571), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n560), .A2(G169), .A3(new_n571), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n560), .A2(KEYINPUT21), .A3(G169), .A4(new_n571), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n569), .A2(new_n573), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n317), .A2(new_n321), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n290), .A2(new_n210), .A3(G68), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n262), .A2(new_n427), .ZN(new_n581));
  XOR2_X1   g0381(.A(KEYINPUT82), .B(G87), .Z(new_n582));
  NOR3_X1   g0382(.A1(new_n582), .A2(G97), .A3(G107), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n287), .A2(new_n427), .ZN(new_n584));
  AOI21_X1  g0384(.A(G20), .B1(new_n584), .B2(KEYINPUT19), .ZN(new_n585));
  OAI221_X1 g0385(.A(new_n580), .B1(KEYINPUT19), .B2(new_n581), .C1(new_n583), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n579), .B1(new_n586), .B2(new_n271), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n543), .A2(new_n321), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n290), .A2(G244), .A3(G1698), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G116), .ZN(new_n590));
  OAI211_X1 g0390(.A(G238), .B(new_n292), .C1(new_n350), .C2(new_n351), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n296), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n493), .A2(G274), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n298), .A2(G250), .A3(new_n502), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n587), .A2(new_n588), .B1(new_n313), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n596), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n345), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(KEYINPUT81), .A3(new_n345), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n462), .A2(new_n354), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n579), .B(new_n604), .C1(new_n586), .C2(new_n271), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n596), .A2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n302), .C2(new_n596), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n479), .A2(new_n271), .ZN(new_n609));
  INV_X1    g0409(.A(new_n463), .ZN(new_n610));
  INV_X1    g0410(.A(new_n465), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n507), .A2(G169), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n506), .A2(new_n485), .A3(KEYINPUT86), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT86), .B1(new_n506), .B2(new_n485), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n499), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n616), .B2(new_n345), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT87), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT87), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n612), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n608), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n461), .A2(new_n551), .A3(new_n578), .A4(new_n622), .ZN(G372));
  OAI21_X1  g0423(.A(KEYINPUT26), .B1(new_n608), .B2(new_n550), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n597), .A2(new_n599), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n607), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n550), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n551), .A2(new_n607), .A3(new_n625), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n576), .A2(new_n569), .A3(new_n577), .ZN(new_n632));
  INV_X1    g0432(.A(new_n618), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n624), .B(new_n630), .C1(new_n631), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n461), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n315), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n389), .A2(new_n405), .A3(new_n407), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT18), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n408), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n348), .A2(new_n457), .B1(new_n441), .B2(new_n453), .ZN(new_n642));
  INV_X1    g0442(.A(new_n401), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n637), .B1(new_n644), .B2(new_n311), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n636), .A2(new_n645), .ZN(G369));
  NOR2_X1   g0446(.A1(new_n273), .A2(G20), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n214), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n560), .A2(new_n653), .ZN(new_n654));
  MUX2_X1   g0454(.A(new_n632), .B(new_n578), .S(new_n654), .Z(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n619), .A2(new_n621), .ZN(new_n657));
  INV_X1    g0457(.A(new_n653), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n515), .C1(new_n480), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n633), .A2(new_n653), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n515), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n632), .A2(new_n658), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n653), .B(KEYINPUT88), .Z(new_n668));
  NOR2_X1   g0468(.A1(new_n618), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n217), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G1), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n583), .A2(new_n224), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n675), .A2(new_n676), .B1(new_n209), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  INV_X1    g0479(.A(new_n668), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n635), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n550), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n629), .A3(new_n607), .A4(new_n603), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n627), .B2(new_n550), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n625), .A2(KEYINPUT92), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n657), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n632), .ZN(new_n688));
  OAI221_X1 g0488(.A(new_n686), .B1(KEYINPUT92), .B2(new_n625), .C1(new_n688), .C2(new_n631), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(new_n658), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n681), .B1(new_n690), .B2(new_n679), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n571), .A2(new_n596), .A3(new_n345), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT90), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n571), .A2(new_n596), .A3(new_n694), .A4(new_n345), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n530), .A3(new_n616), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT89), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n596), .B1(new_n511), .B2(new_n512), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n547), .A2(new_n567), .ZN(new_n701));
  AOI211_X1 g0501(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n513), .A2(new_n532), .A3(new_n568), .A4(new_n598), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT30), .B1(new_n703), .B2(KEYINPUT89), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n697), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT91), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n697), .B(KEYINPUT91), .C1(new_n702), .C2(new_n704), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n653), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n622), .A2(new_n578), .A3(new_n551), .A4(new_n680), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n691), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n678), .B1(new_n717), .B2(G1), .ZN(G364));
  AOI21_X1  g0518(.A(new_n675), .B1(G45), .B2(new_n647), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n655), .B2(G330), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G330), .B2(new_n655), .ZN(new_n721));
  INV_X1    g0521(.A(new_n719), .ZN(new_n722));
  NOR4_X1   g0522(.A1(new_n210), .A2(new_n302), .A3(new_n365), .A4(G179), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n210), .A2(new_n345), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(new_n302), .A3(G200), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G322), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n371), .B1(new_n563), .B2(new_n724), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n725), .A2(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G190), .ZN(new_n732));
  INV_X1    g0532(.A(G317), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT33), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(KEYINPUT33), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G283), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n210), .A2(G190), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n345), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n302), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n210), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n736), .B1(new_n737), .B2(new_n739), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n730), .B(new_n743), .C1(G311), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n731), .A2(new_n302), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G326), .ZN(new_n747));
  INV_X1    g0547(.A(G329), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n738), .A2(new_n345), .A3(new_n365), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT93), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n745), .B(new_n747), .C1(new_n748), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n739), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G107), .ZN(new_n760));
  INV_X1    g0560(.A(new_n746), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n761), .B2(new_n272), .ZN(new_n762));
  INV_X1    g0562(.A(new_n267), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n371), .B1(new_n727), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n723), .A2(new_n582), .ZN(new_n765));
  INV_X1    g0565(.A(new_n744), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n764), .B(new_n765), .C1(new_n253), .C2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n762), .B(new_n767), .C1(G68), .C2(new_n732), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  OR3_X1    g0569(.A1(new_n753), .A2(KEYINPUT32), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(KEYINPUT32), .B1(new_n753), .B2(new_n769), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n742), .A2(new_n427), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n758), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n211), .B1(G20), .B2(new_n313), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n775), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n672), .A2(new_n290), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n206), .A2(new_n492), .A3(G50), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n780), .B(new_n781), .C1(new_n254), .C2(new_n492), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n672), .A2(new_n371), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G355), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n782), .B(new_n784), .C1(G116), .C2(new_n217), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n774), .A2(new_n775), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n778), .B(KEYINPUT95), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n655), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n721), .B1(new_n722), .B2(new_n789), .ZN(G396));
  AOI22_X1  g0590(.A1(G116), .A2(new_n744), .B1(new_n732), .B2(G283), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT96), .Z(new_n792));
  AOI211_X1 g0592(.A(new_n773), .B(new_n792), .C1(G303), .C2(new_n746), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n371), .B1(new_n336), .B2(new_n724), .C1(new_n728), .C2(new_n740), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G87), .B2(new_n759), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n793), .B(new_n795), .C1(new_n796), .C2(new_n757), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n739), .A2(new_n202), .ZN(new_n798));
  INV_X1    g0598(.A(new_n742), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n763), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n727), .A2(G143), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n744), .A2(G159), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n732), .A2(G150), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n746), .A2(G137), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n290), .B1(new_n724), .B2(new_n272), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n805), .B2(new_n806), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n757), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n797), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n775), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n775), .A2(new_n776), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n333), .A2(new_n653), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n348), .B1(new_n425), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n347), .A2(new_n653), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n813), .B1(G77), .B2(new_n815), .C1(new_n819), .C2(new_n777), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n719), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n635), .A2(new_n680), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(new_n819), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(new_n715), .Z(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n824), .B2(new_n719), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT97), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  NAND3_X1  g0627(.A1(new_n441), .A2(new_n453), .A3(new_n658), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT39), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n394), .A2(new_n398), .A3(new_n388), .ZN(new_n830));
  INV_X1    g0630(.A(new_n651), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n389), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n638), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n638), .A2(new_n830), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(KEYINPUT98), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n834), .A2(new_n836), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n832), .B1(new_n641), .B2(new_n401), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT38), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n832), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n410), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n838), .A3(new_n837), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n840), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AND4_X1   g0647(.A1(KEYINPUT98), .A2(new_n842), .A3(new_n838), .A4(new_n837), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n829), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n843), .A2(KEYINPUT39), .A3(new_n846), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n828), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n818), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n822), .B2(new_n817), .ZN(new_n853));
  INV_X1    g0653(.A(new_n457), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n453), .B(new_n653), .C1(new_n854), .C2(new_n441), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n454), .B(new_n457), .C1(new_n452), .C2(new_n658), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND4_X1   g0657(.A1(new_n843), .A2(new_n853), .A3(new_n846), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n641), .A2(new_n831), .ZN(new_n859));
  OR3_X1    g0659(.A1(new_n851), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n461), .A2(new_n691), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n861), .A2(new_n645), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n860), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n711), .A2(KEYINPUT99), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n653), .A4(new_n708), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(new_n712), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT99), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n709), .A2(new_n867), .A3(new_n710), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n425), .A2(new_n816), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n347), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n857), .A2(new_n871), .A3(new_n852), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT100), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT38), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n838), .B1(new_n845), .B2(new_n837), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n839), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n848), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT40), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n874), .B2(new_n875), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT100), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT40), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n869), .A3(new_n872), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n461), .A2(new_n869), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(G330), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n863), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n214), .B2(new_n647), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n224), .B1(new_n539), .B2(KEYINPUT35), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n211), .A2(new_n210), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n891), .B(new_n892), .C1(KEYINPUT35), .C2(new_n539), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT36), .ZN(new_n894));
  OAI21_X1  g0694(.A(G77), .B1(new_n267), .B2(new_n202), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n209), .A2(new_n895), .B1(G50), .B2(new_n202), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n273), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT101), .Z(G367));
  NOR2_X1   g0699(.A1(new_n739), .A2(new_n253), .ZN(new_n900));
  INV_X1    g0700(.A(G137), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n290), .B1(new_n267), .B2(new_n724), .C1(new_n753), .C2(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n900), .B(new_n902), .C1(G143), .C2(new_n746), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G50), .A2(new_n744), .B1(new_n732), .B2(G159), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT108), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n742), .A2(new_n202), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(G150), .B2(new_n727), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n903), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT109), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT46), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n724), .B2(new_n224), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n759), .A2(G97), .ZN(new_n913));
  INV_X1    g0713(.A(new_n732), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n912), .B(new_n913), .C1(new_n740), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(G311), .B2(new_n746), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n724), .A2(new_n911), .A3(new_n224), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(G107), .B2(new_n799), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n290), .B1(new_n727), .B2(G303), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n920), .B1(new_n737), .B2(new_n766), .C1(new_n733), .C2(new_n753), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT47), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n775), .ZN(new_n924));
  INV_X1    g0724(.A(new_n780), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n779), .B1(new_n217), .B2(new_n322), .C1(new_n245), .C2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT102), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n605), .A2(new_n658), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n627), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n626), .A2(new_n928), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT102), .B1(new_n626), .B2(new_n928), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n787), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n924), .A2(new_n719), .A3(new_n926), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n214), .B1(new_n647), .B2(G45), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n682), .A2(new_n668), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n546), .A2(new_n668), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n545), .A2(new_n550), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n670), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT45), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT44), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT104), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n667), .A2(new_n669), .ZN(new_n947));
  INV_X1    g0747(.A(new_n941), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n670), .A2(KEYINPUT104), .A3(new_n941), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n946), .A3(new_n948), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT104), .B1(new_n670), .B2(new_n941), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(KEYINPUT44), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n944), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n937), .B1(new_n955), .B2(new_n663), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n663), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n944), .A2(new_n951), .A3(new_n664), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n956), .B1(new_n959), .B2(new_n937), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n662), .A2(new_n666), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n665), .B2(new_n666), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n656), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n716), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n716), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n673), .B(KEYINPUT41), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n936), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT106), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n667), .A2(new_n941), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n970), .A2(KEYINPUT103), .A3(KEYINPUT42), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(KEYINPUT42), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT103), .B1(new_n970), .B2(KEYINPUT42), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n687), .A2(new_n545), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n680), .B1(new_n974), .B2(new_n682), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT43), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(new_n933), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n663), .A2(new_n941), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n933), .A2(new_n977), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n968), .A2(new_n969), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n969), .B1(new_n968), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n935), .B1(new_n984), .B2(new_n985), .ZN(G387));
  INV_X1    g0786(.A(new_n964), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n673), .B(KEYINPUT114), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n716), .A2(new_n963), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n242), .A2(new_n492), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n992), .A2(new_n780), .B1(new_n676), .B2(new_n783), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n320), .A2(G50), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT50), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n202), .B2(new_n253), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n996), .A2(G45), .A3(new_n676), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n993), .A2(new_n997), .B1(G107), .B2(new_n217), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n722), .B1(new_n998), .B2(new_n779), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  AND2_X1   g0800(.A1(new_n754), .A2(G326), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n744), .A2(G303), .B1(new_n746), .B2(G322), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n796), .B2(new_n914), .C1(new_n733), .C2(new_n728), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n1005));
  AOI22_X1  g0805(.A1(new_n1004), .A2(new_n1005), .B1(G283), .B2(new_n799), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n740), .B2(new_n724), .C1(new_n1005), .C2(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n290), .B(new_n1001), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .C1(new_n224), .C2(new_n739), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n913), .B1(new_n753), .B2(new_n257), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n322), .A2(new_n742), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n290), .B1(new_n253), .B2(new_n724), .C1(new_n728), .C2(new_n272), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G159), .C2(new_n746), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n766), .A2(new_n202), .B1(new_n914), .B2(new_n268), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT111), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1010), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n775), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1000), .B1(new_n661), .B2(new_n788), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n991), .B(new_n1021), .C1(new_n936), .C2(new_n963), .ZN(G393));
  NAND2_X1  g0822(.A1(new_n960), .A2(new_n964), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n988), .B1(new_n987), .B2(new_n959), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n936), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n957), .A2(new_n1026), .A3(new_n958), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n727), .A2(G159), .B1(new_n746), .B2(G150), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT51), .Z(new_n1029));
  OAI221_X1 g0829(.A(new_n290), .B1(new_n202), .B2(new_n724), .C1(new_n766), .C2(new_n320), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G77), .B2(new_n799), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n754), .A2(G143), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n732), .A2(G50), .B1(new_n759), .B2(G87), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n290), .B1(new_n723), .B2(G283), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n760), .B(new_n1035), .C1(new_n753), .C2(new_n729), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT115), .Z(new_n1037));
  AOI22_X1  g0837(.A1(new_n727), .A2(G311), .B1(new_n746), .B2(G317), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT52), .Z(new_n1039));
  AOI22_X1  g0839(.A1(G116), .A2(new_n799), .B1(new_n732), .B2(G303), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n766), .A2(new_n740), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n722), .B1(new_n1043), .B2(new_n775), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n779), .B1(new_n427), .B2(new_n217), .C1(new_n250), .C2(new_n925), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n778), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1044), .B(new_n1045), .C1(new_n1046), .C2(new_n941), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1025), .A2(new_n1027), .A3(new_n1047), .ZN(G390));
  NAND2_X1  g0848(.A1(new_n853), .A2(new_n857), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n828), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n849), .A3(new_n850), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n689), .A2(new_n658), .A3(new_n871), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n852), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n857), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n847), .A2(new_n848), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n828), .A3(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n714), .A2(G330), .A3(new_n819), .A4(new_n857), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1051), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n869), .A2(G330), .A3(new_n819), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n857), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n459), .A2(new_n460), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n459), .A2(new_n460), .ZN(new_n1066));
  OAI211_X1 g0866(.A(G330), .B(new_n869), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n861), .A2(new_n645), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(G330), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n817), .A2(new_n1069), .A3(new_n818), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n857), .B1(new_n1070), .B2(new_n714), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n853), .B1(new_n1062), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1053), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT116), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1060), .A2(new_n1061), .B1(KEYINPUT116), .B2(new_n1057), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1068), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1064), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1068), .B(new_n1078), .C1(new_n1059), .C2(new_n1063), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n989), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1026), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n849), .A2(new_n776), .A3(new_n850), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n728), .A2(new_n224), .B1(new_n253), .B2(new_n742), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT117), .Z(new_n1086));
  OAI221_X1 g0886(.A(new_n371), .B1(new_n354), .B2(new_n724), .C1(new_n766), .C2(new_n427), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n914), .A2(new_n336), .ZN(new_n1088));
  NOR4_X1   g0888(.A1(new_n1086), .A2(new_n798), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n737), .B2(new_n761), .C1(new_n740), .C2(new_n757), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n732), .A2(G137), .B1(new_n759), .B2(G50), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n761), .C1(new_n769), .C2(new_n742), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n723), .A2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n290), .B1(new_n728), .B2(new_n810), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  INV_X1    g0898(.A(G125), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1097), .B1(new_n766), .B2(new_n1098), .C1(new_n1099), .C2(new_n757), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1020), .B1(new_n1090), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n268), .B2(new_n814), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1084), .A2(new_n719), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1082), .A2(new_n1083), .A3(new_n1103), .ZN(G378));
  INV_X1    g0904(.A(KEYINPUT57), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1081), .B2(new_n1068), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n851), .A2(new_n858), .A3(new_n859), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT56), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT55), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n282), .A2(new_n651), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n316), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1110), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n311), .A2(new_n315), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1109), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1112), .B1(new_n311), .B2(new_n315), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n637), .B(new_n1110), .C1(new_n308), .C2(new_n310), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT55), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1111), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT55), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(KEYINPUT56), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n885), .B2(G330), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1069), .B(new_n1122), .C1(new_n879), .C2(new_n884), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1107), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n884), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n709), .A2(new_n867), .A3(new_n710), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n867), .B1(new_n709), .B2(new_n710), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n865), .A2(new_n712), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n819), .A2(new_n857), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n882), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1055), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1127), .B1(new_n1134), .B2(KEYINPUT40), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1122), .B1(new_n1135), .B2(new_n1069), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n885), .A2(G330), .A3(new_n1123), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n860), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT121), .B1(new_n1126), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n860), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT121), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1106), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT120), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1124), .A2(new_n1125), .A3(new_n1107), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n1140), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1126), .A2(new_n1138), .A3(KEYINPUT120), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1146), .A2(new_n1147), .B1(new_n1068), .B2(new_n1081), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n989), .B(new_n1143), .C1(new_n1148), .C2(KEYINPUT57), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1123), .A2(new_n776), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n488), .B1(new_n253), .B2(new_n724), .C1(new_n757), .C2(new_n737), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n739), .A2(new_n267), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n290), .A3(new_n1152), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT118), .Z(new_n1154));
  OAI22_X1  g0954(.A1(new_n914), .A2(new_n427), .B1(new_n761), .B2(new_n224), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n906), .B(new_n1155), .C1(new_n321), .C2(new_n744), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(new_n336), .C2(new_n728), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT58), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n914), .A2(new_n810), .B1(new_n761), .B2(new_n1099), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G128), .A2(new_n727), .B1(new_n744), .B2(G137), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n724), .B2(new_n1098), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G150), .C2(new_n799), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n754), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G33), .B1(new_n759), .B2(G159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n272), .B1(new_n350), .B2(G41), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1159), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n775), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n719), .B1(G50), .B2(new_n815), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT119), .Z(new_n1173));
  NAND3_X1  g0973(.A1(new_n1150), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n1026), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1149), .A2(new_n1177), .ZN(G375));
  OR2_X1    g0978(.A1(new_n1068), .A2(new_n1078), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n966), .A3(new_n1079), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n728), .A2(new_n901), .B1(new_n914), .B2(new_n1098), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n290), .B1(new_n766), .B2(new_n257), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1152), .B(new_n1182), .C1(G50), .C2(new_n799), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n769), .B2(new_n724), .C1(new_n757), .C2(new_n1092), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT124), .Z(new_n1185));
  AOI211_X1 g0985(.A(new_n1181), .B(new_n1185), .C1(G132), .C2(new_n746), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n371), .B1(new_n766), .B2(new_n336), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G97), .B2(new_n723), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n727), .A2(G283), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1012), .A2(new_n900), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n746), .A2(G294), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n757), .A2(new_n563), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G116), .C2(new_n732), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1186), .A2(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1195), .A2(new_n1020), .B1(new_n777), .B2(new_n857), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n719), .B1(G68), .B2(new_n815), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT123), .Z(new_n1198));
  NOR2_X1   g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n936), .B(KEYINPUT122), .Z(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1078), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1180), .A2(new_n1201), .ZN(G381));
  INV_X1    g1002(.A(G378), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1149), .A2(new_n1203), .A3(new_n1177), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1204), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n935), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n968), .A2(new_n982), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT106), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n1208), .B2(new_n983), .ZN(new_n1209));
  INV_X1    g1009(.A(G390), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n826), .A3(new_n1209), .A4(new_n1210), .ZN(G407));
  OAI211_X1 g1011(.A(G407), .B(G213), .C1(G343), .C2(new_n1204), .ZN(G409));
  INV_X1    g1012(.A(KEYINPUT126), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT63), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1081), .A2(new_n1068), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1143), .A2(new_n989), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G378), .B(new_n1177), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT125), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT125), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1149), .A2(new_n1220), .A3(G378), .A4(new_n1177), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1200), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1126), .A2(new_n1138), .A3(KEYINPUT120), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT120), .B1(new_n1126), .B2(new_n1138), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1215), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1174), .B(new_n1223), .C1(new_n1226), .C2(new_n967), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n1203), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1222), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G343), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n988), .B1(new_n1179), .B2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1235), .B(new_n1079), .C1(new_n1234), .C2(new_n1179), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n826), .A3(new_n1201), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n826), .B1(new_n1236), .B2(new_n1201), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1230), .A2(new_n1233), .A3(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G2897), .B(new_n1232), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1239), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1232), .A2(G2897), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1237), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1228), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n1232), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1214), .B1(new_n1242), .B2(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(G393), .B(G396), .Z(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1208), .A2(new_n983), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G390), .B1(new_n1253), .B2(new_n935), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1206), .B(new_n1210), .C1(new_n1208), .C2(new_n983), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1210), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1209), .A2(G390), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1251), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1256), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1248), .A2(new_n1232), .A3(new_n1240), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(KEYINPUT63), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1213), .B1(new_n1250), .B2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT63), .B1(new_n1266), .B2(new_n1262), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1256), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1242), .B2(new_n1214), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(KEYINPUT126), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1232), .B1(new_n1222), .B2(new_n1229), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT127), .B1(new_n1273), .B2(new_n1241), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT127), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1248), .A2(new_n1275), .A3(new_n1232), .A4(new_n1240), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1274), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1273), .A2(KEYINPUT127), .A3(new_n1241), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1260), .B(new_n1249), .C1(new_n1279), .C2(KEYINPUT62), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1272), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1271), .A2(new_n1281), .ZN(G405));
  XNOR2_X1  g1082(.A(new_n1272), .B(new_n1240), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1219), .A2(new_n1221), .B1(new_n1203), .B2(G375), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1283), .B(new_n1284), .ZN(G402));
endmodule


