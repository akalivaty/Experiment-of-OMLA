

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U323 ( .A(n414), .B(n413), .ZN(n422) );
  XNOR2_X1 U324 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n413) );
  XNOR2_X1 U325 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U326 ( .A(n406), .B(n405), .ZN(n409) );
  XNOR2_X1 U327 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U328 ( .A(n424), .B(n423), .ZN(n552) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n423) );
  NOR2_X1 U330 ( .A1(n422), .A2(n421), .ZN(n424) );
  NOR2_X1 U331 ( .A1(n468), .A2(n420), .ZN(n421) );
  XNOR2_X1 U332 ( .A(n387), .B(n342), .ZN(n343) );
  XNOR2_X1 U333 ( .A(n386), .B(n385), .ZN(n391) );
  XOR2_X1 U334 ( .A(n411), .B(n410), .Z(n567) );
  INV_X1 U335 ( .A(n552), .ZN(n553) );
  XOR2_X1 U336 ( .A(G134GAT), .B(G106GAT), .Z(n291) );
  XNOR2_X1 U337 ( .A(n341), .B(KEYINPUT15), .ZN(n342) );
  INV_X1 U338 ( .A(KEYINPUT32), .ZN(n375) );
  INV_X1 U339 ( .A(KEYINPUT54), .ZN(n435) );
  INV_X1 U340 ( .A(n398), .ZN(n399) );
  XNOR2_X1 U341 ( .A(n435), .B(KEYINPUT119), .ZN(n436) );
  INV_X1 U342 ( .A(KEYINPUT77), .ZN(n403) );
  XNOR2_X1 U343 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U344 ( .A(n349), .B(n348), .ZN(n350) );
  NOR2_X1 U345 ( .A1(n481), .A2(n579), .ZN(n460) );
  XNOR2_X1 U346 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U347 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U348 ( .A(n407), .B(n291), .ZN(n408) );
  XNOR2_X1 U349 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U350 ( .A(n462), .B(KEYINPUT120), .ZN(n576) );
  XOR2_X1 U351 ( .A(n481), .B(KEYINPUT28), .Z(n533) );
  XNOR2_X1 U352 ( .A(n465), .B(G190GAT), .ZN(n466) );
  XNOR2_X1 U353 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XOR2_X1 U354 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n293) );
  XNOR2_X1 U355 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n292) );
  XNOR2_X1 U356 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U357 ( .A(G169GAT), .B(n294), .Z(n432) );
  XOR2_X1 U358 ( .A(KEYINPUT0), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U359 ( .A(KEYINPUT83), .B(G120GAT), .ZN(n295) );
  XNOR2_X1 U360 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U361 ( .A(G113GAT), .B(n297), .Z(n454) );
  XNOR2_X1 U362 ( .A(n432), .B(n454), .ZN(n310) );
  XOR2_X1 U363 ( .A(KEYINPUT20), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U365 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U366 ( .A(G71GAT), .B(KEYINPUT86), .Z(n301) );
  XNOR2_X1 U367 ( .A(KEYINPUT65), .B(KEYINPUT84), .ZN(n300) );
  XNOR2_X1 U368 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U369 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G127GAT), .Z(n345) );
  XOR2_X1 U371 ( .A(G183GAT), .B(G176GAT), .Z(n305) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U373 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U374 ( .A(n345), .B(n306), .ZN(n307) );
  XNOR2_X1 U375 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U376 ( .A(n310), .B(n309), .ZN(n536) );
  XOR2_X1 U377 ( .A(KEYINPUT24), .B(G218GAT), .Z(n312) );
  XOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT21), .Z(n425) );
  XOR2_X1 U379 ( .A(G22GAT), .B(G155GAT), .Z(n344) );
  XNOR2_X1 U380 ( .A(n425), .B(n344), .ZN(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U382 ( .A(G50GAT), .B(G162GAT), .Z(n398) );
  XOR2_X1 U383 ( .A(n313), .B(n398), .Z(n318) );
  XOR2_X1 U384 ( .A(KEYINPUT22), .B(G204GAT), .Z(n315) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U386 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U387 ( .A(KEYINPUT88), .B(n316), .ZN(n317) );
  XNOR2_X1 U388 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U389 ( .A(KEYINPUT23), .B(G211GAT), .Z(n320) );
  XNOR2_X1 U390 ( .A(KEYINPUT87), .B(KEYINPUT89), .ZN(n319) );
  XNOR2_X1 U391 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U392 ( .A(n322), .B(n321), .Z(n331) );
  INV_X1 U393 ( .A(G148GAT), .ZN(n323) );
  NAND2_X1 U394 ( .A1(G78GAT), .A2(n323), .ZN(n326) );
  INV_X1 U395 ( .A(G78GAT), .ZN(n324) );
  NAND2_X1 U396 ( .A1(n324), .A2(G148GAT), .ZN(n325) );
  NAND2_X1 U397 ( .A1(n326), .A2(n325), .ZN(n328) );
  XNOR2_X1 U398 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n327) );
  XNOR2_X1 U399 ( .A(n328), .B(n327), .ZN(n378) );
  XNOR2_X1 U400 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n329) );
  XNOR2_X1 U401 ( .A(n329), .B(KEYINPUT2), .ZN(n450) );
  XNOR2_X1 U402 ( .A(n378), .B(n450), .ZN(n330) );
  XNOR2_X1 U403 ( .A(n331), .B(n330), .ZN(n481) );
  XOR2_X1 U404 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n333) );
  XNOR2_X1 U405 ( .A(KEYINPUT80), .B(KEYINPUT12), .ZN(n332) );
  XNOR2_X1 U406 ( .A(n333), .B(n332), .ZN(n353) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U408 ( .A(n334), .B(G211GAT), .ZN(n429) );
  INV_X1 U409 ( .A(KEYINPUT13), .ZN(n335) );
  NAND2_X1 U410 ( .A1(G57GAT), .A2(n335), .ZN(n338) );
  INV_X1 U411 ( .A(G57GAT), .ZN(n336) );
  NAND2_X1 U412 ( .A1(n336), .A2(KEYINPUT13), .ZN(n337) );
  NAND2_X1 U413 ( .A1(n338), .A2(n337), .ZN(n340) );
  XNOR2_X1 U414 ( .A(G71GAT), .B(KEYINPUT72), .ZN(n339) );
  XNOR2_X1 U415 ( .A(n340), .B(n339), .ZN(n387) );
  AND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XOR2_X1 U417 ( .A(n429), .B(n343), .Z(n347) );
  XNOR2_X1 U418 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U419 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U420 ( .A(KEYINPUT71), .B(G1GAT), .Z(n366) );
  XNOR2_X1 U421 ( .A(n366), .B(G78GAT), .ZN(n349) );
  INV_X1 U422 ( .A(G64GAT), .ZN(n348) );
  XOR2_X1 U423 ( .A(n353), .B(n352), .Z(n415) );
  XOR2_X1 U424 ( .A(KEYINPUT109), .B(n415), .Z(n575) );
  XOR2_X1 U425 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n355) );
  XNOR2_X1 U426 ( .A(G8GAT), .B(KEYINPUT66), .ZN(n354) );
  XNOR2_X1 U427 ( .A(n355), .B(n354), .ZN(n374) );
  XOR2_X1 U428 ( .A(G22GAT), .B(G197GAT), .Z(n357) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(G50GAT), .ZN(n356) );
  XNOR2_X1 U430 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U431 ( .A(G113GAT), .B(G15GAT), .Z(n359) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U433 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U434 ( .A(n361), .B(n360), .Z(n372) );
  XOR2_X1 U435 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n363) );
  XNOR2_X1 U436 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n362) );
  XNOR2_X1 U437 ( .A(n363), .B(n362), .ZN(n370) );
  XOR2_X1 U438 ( .A(G29GAT), .B(G43GAT), .Z(n365) );
  XNOR2_X1 U439 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n364) );
  XNOR2_X1 U440 ( .A(n365), .B(n364), .ZN(n402) );
  XOR2_X1 U441 ( .A(n402), .B(n366), .Z(n368) );
  NAND2_X1 U442 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U443 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U444 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U445 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n374), .B(n373), .ZN(n581) );
  INV_X1 U447 ( .A(n581), .ZN(n555) );
  NAND2_X1 U448 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  INV_X1 U449 ( .A(KEYINPUT33), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n386) );
  XOR2_X1 U451 ( .A(G99GAT), .B(G85GAT), .Z(n407) );
  XNOR2_X1 U452 ( .A(G120GAT), .B(n407), .ZN(n384) );
  XOR2_X1 U453 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n382) );
  XNOR2_X1 U454 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U456 ( .A(G64GAT), .B(G92GAT), .Z(n389) );
  XNOR2_X1 U457 ( .A(G176GAT), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n426) );
  XOR2_X1 U459 ( .A(n387), .B(n426), .Z(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n468) );
  XNOR2_X1 U461 ( .A(KEYINPUT41), .B(n468), .ZN(n571) );
  NOR2_X1 U462 ( .A1(n555), .A2(n571), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n392), .B(KEYINPUT46), .ZN(n393) );
  NOR2_X1 U464 ( .A1(n575), .A2(n393), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n394), .B(KEYINPUT110), .ZN(n412) );
  XOR2_X1 U466 ( .A(KEYINPUT10), .B(G92GAT), .Z(n396) );
  XNOR2_X1 U467 ( .A(KEYINPUT78), .B(KEYINPUT11), .ZN(n395) );
  XNOR2_X1 U468 ( .A(n396), .B(n395), .ZN(n411) );
  XNOR2_X1 U469 ( .A(G36GAT), .B(G190GAT), .ZN(n397) );
  XNOR2_X1 U470 ( .A(n397), .B(G218GAT), .ZN(n431) );
  XNOR2_X1 U471 ( .A(n431), .B(n399), .ZN(n401) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U473 ( .A(n401), .B(n400), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n402), .B(KEYINPUT9), .ZN(n404) );
  AND2_X1 U475 ( .A1(n412), .A2(n567), .ZN(n414) );
  XNOR2_X1 U476 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n416) );
  XOR2_X1 U477 ( .A(n416), .B(n567), .Z(n589) );
  NAND2_X1 U478 ( .A1(n415), .A2(n589), .ZN(n418) );
  XOR2_X1 U479 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U481 ( .A1(n419), .A2(n555), .ZN(n420) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U483 ( .A1(G226GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n526) );
  NOR2_X1 U488 ( .A1(n552), .A2(n526), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n459) );
  XOR2_X1 U490 ( .A(G57GAT), .B(G148GAT), .Z(n439) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(G127GAT), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U493 ( .A(G85GAT), .B(G155GAT), .Z(n441) );
  XNOR2_X1 U494 ( .A(G29GAT), .B(G162GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n458) );
  XOR2_X1 U497 ( .A(KEYINPUT4), .B(KEYINPUT94), .Z(n445) );
  XNOR2_X1 U498 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n447) );
  XNOR2_X1 U501 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n456) );
  XOR2_X1 U504 ( .A(n450), .B(KEYINPUT1), .Z(n452) );
  NAND2_X1 U505 ( .A1(G225GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U509 ( .A(n458), .B(n457), .Z(n477) );
  INV_X1 U510 ( .A(n477), .ZN(n524) );
  NAND2_X1 U511 ( .A1(n459), .A2(n524), .ZN(n579) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT55), .ZN(n461) );
  NOR2_X1 U513 ( .A1(n536), .A2(n461), .ZN(n462) );
  AND2_X1 U514 ( .A1(n576), .A2(n581), .ZN(n464) );
  XNOR2_X1 U515 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n464), .B(n463), .ZN(G1348GAT) );
  INV_X1 U517 ( .A(n567), .ZN(n547) );
  NAND2_X1 U518 ( .A1(n576), .A2(n547), .ZN(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n465) );
  NOR2_X1 U520 ( .A1(n555), .A2(n468), .ZN(n501) );
  NOR2_X1 U521 ( .A1(n536), .A2(n526), .ZN(n469) );
  XOR2_X1 U522 ( .A(KEYINPUT97), .B(n469), .Z(n470) );
  NOR2_X1 U523 ( .A1(n481), .A2(n470), .ZN(n471) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n471), .Z(n475) );
  XNOR2_X1 U525 ( .A(n526), .B(KEYINPUT27), .ZN(n479) );
  NAND2_X1 U526 ( .A1(n481), .A2(n536), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT96), .ZN(n473) );
  XNOR2_X1 U528 ( .A(KEYINPUT26), .B(n473), .ZN(n578) );
  NOR2_X1 U529 ( .A1(n479), .A2(n578), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(n478), .Z(n484) );
  NOR2_X1 U533 ( .A1(n479), .A2(n524), .ZN(n480) );
  XNOR2_X1 U534 ( .A(n480), .B(KEYINPUT95), .ZN(n551) );
  INV_X1 U535 ( .A(n533), .ZN(n482) );
  NOR2_X1 U536 ( .A1(n551), .A2(n482), .ZN(n538) );
  NAND2_X1 U537 ( .A1(n536), .A2(n538), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n484), .A2(n483), .ZN(n498) );
  XOR2_X1 U539 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n486) );
  NAND2_X1 U540 ( .A1(n415), .A2(n567), .ZN(n485) );
  XNOR2_X1 U541 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  AND2_X1 U543 ( .A1(n498), .A2(n488), .ZN(n514) );
  NAND2_X1 U544 ( .A1(n501), .A2(n514), .ZN(n496) );
  NOR2_X1 U545 ( .A1(n524), .A2(n496), .ZN(n489) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(n489), .Z(n490) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U548 ( .A1(n526), .A2(n496), .ZN(n492) );
  XNOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n493), .ZN(G1325GAT) );
  NOR2_X1 U552 ( .A1(n536), .A2(n496), .ZN(n495) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U555 ( .A1(n533), .A2(n496), .ZN(n497) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NAND2_X1 U557 ( .A1(n589), .A2(n498), .ZN(n499) );
  NOR2_X1 U558 ( .A1(n415), .A2(n499), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT37), .B(n500), .Z(n523) );
  NAND2_X1 U560 ( .A1(n523), .A2(n501), .ZN(n503) );
  XOR2_X1 U561 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(n511) );
  NOR2_X1 U563 ( .A1(n511), .A2(n524), .ZN(n507) );
  XOR2_X1 U564 ( .A(KEYINPUT101), .B(KEYINPUT104), .Z(n505) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n526), .A2(n511), .ZN(n508) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n508), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n536), .A2(n511), .ZN(n509) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(n509), .Z(n510) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n513) );
  NOR2_X1 U574 ( .A1(n533), .A2(n511), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  NOR2_X1 U576 ( .A1(n581), .A2(n571), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n522), .A2(n514), .ZN(n519) );
  NOR2_X1 U578 ( .A1(n524), .A2(n519), .ZN(n515) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n519), .ZN(n517) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n536), .A2(n519), .ZN(n518) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n518), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n533), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n532) );
  NOR2_X1 U589 ( .A1(n524), .A2(n532), .ZN(n525) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n532), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT106), .B(n527), .Z(n528) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NOR2_X1 U594 ( .A1(n536), .A2(n532), .ZN(n529) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT108), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(n535), .B(n534), .Z(G1339GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n552), .ZN(n537) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U603 ( .A1(n555), .A2(n544), .ZN(n539) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U605 ( .A1(n544), .A2(n571), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n541) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT113), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  INV_X1 U610 ( .A(n544), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n548), .A2(n575), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n578), .A2(n551), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n566) );
  NOR2_X1 U619 ( .A1(n555), .A2(n566), .ZN(n557) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n559) );
  XNOR2_X1 U623 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n563) );
  NOR2_X1 U625 ( .A1(n566), .A2(n571), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  INV_X1 U629 ( .A(n415), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n564), .A2(n566), .ZN(n565) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n565), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n568), .Z(G1347GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n574) );
  INV_X1 U637 ( .A(n571), .ZN(n572) );
  AND2_X1 U638 ( .A1(n576), .A2(n572), .ZN(n573) );
  XOR2_X1 U639 ( .A(n574), .B(n573), .Z(G1349GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT124), .B(n580), .ZN(n590) );
  AND2_X1 U644 ( .A1(n581), .A2(n590), .ZN(n584) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U649 ( .A1(n468), .A2(n590), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT125), .Z(n588) );
  NAND2_X1 U652 ( .A1(n415), .A2(n590), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n594) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(G1355GAT) );
endmodule

