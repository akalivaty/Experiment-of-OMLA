//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT69), .ZN(new_n203));
  XOR2_X1   g002(.A(G71gat), .B(G99gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT70), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n203), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g013(.A(KEYINPUT1), .B(G127gat), .C1(new_n209), .C2(new_n211), .ZN(new_n215));
  OAI21_X1  g014(.A(G134gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n207), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g018(.A(G127gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n213), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G134gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT25), .B(new_n226), .C1(new_n228), .C2(new_n225), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT24), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n233), .A2(KEYINPUT65), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n230), .A2(new_n239), .A3(new_n231), .A4(new_n232), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n229), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n242), .B1(new_n235), .B2(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n227), .A2(G169gat), .A3(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n225), .ZN(new_n246));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT23), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT25), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT26), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(new_n225), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n234), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(new_n231), .B2(KEYINPUT27), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(new_n230), .A3(new_n232), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT27), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G183gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n231), .A2(KEYINPUT27), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n257), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n231), .A2(KEYINPUT27), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n261), .A2(G183gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT67), .ZN(new_n270));
  AND2_X1   g069(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n271), .A2(new_n272), .A3(new_n257), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n256), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n224), .B1(new_n251), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n233), .A2(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n235), .A2(new_n237), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n240), .ZN(new_n279));
  INV_X1    g078(.A(new_n229), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n226), .B1(new_n228), .B2(new_n225), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n243), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n275), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n222), .B1(new_n219), .B2(new_n221), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G227gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n206), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n294), .B(KEYINPUT32), .C1(new_n295), .C2(new_n206), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n293), .B1(new_n276), .B2(new_n290), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT34), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI211_X1 g102(.A(KEYINPUT34), .B(new_n293), .C1(new_n276), .C2(new_n290), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n298), .A3(new_n299), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT36), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n305), .A2(new_n298), .A3(new_n312), .A4(new_n299), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n307), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT36), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  AND2_X1   g119(.A1(G211gat), .A2(G218gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G211gat), .A2(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G204gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G197gat), .ZN(new_n329));
  INV_X1    g128(.A(G197gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G204gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G211gat), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT73), .A3(new_n325), .ZN(new_n337));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n327), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n320), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT2), .ZN(new_n343));
  INV_X1    g142(.A(G141gat), .ZN(new_n344));
  INV_X1    g143(.A(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G155gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(new_n342), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n342), .ZN(new_n354));
  AND2_X1   g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n354), .B1(new_n357), .B2(new_n343), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n349), .A3(new_n350), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT79), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n348), .A2(new_n362), .A3(KEYINPUT79), .A4(new_n342), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n353), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n341), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n362), .A3(new_n342), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n352), .B1(new_n371), .B2(new_n364), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n333), .A2(new_n339), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT3), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT82), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G228gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(new_n292), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n368), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n320), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n373), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT83), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n341), .A2(new_n366), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(KEYINPUT82), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT3), .B(new_n352), .C1(new_n371), .C2(new_n364), .ZN(new_n388));
  INV_X1    g187(.A(new_n381), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n340), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n386), .A2(new_n387), .A3(new_n390), .A4(new_n368), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n321), .A2(new_n322), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n332), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n381), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n372), .B1(new_n320), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n384), .B1(new_n382), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n383), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G22gat), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n391), .A3(new_n399), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT84), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n406), .A3(new_n400), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n405), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n398), .A2(new_n406), .A3(new_n400), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n372), .A2(new_n224), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n366), .A2(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n380), .A3(new_n289), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n372), .A2(new_n224), .A3(KEYINPUT4), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n366), .A2(new_n289), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n414), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n372), .A2(new_n224), .A3(new_n415), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n372), .A2(new_n224), .A3(KEYINPUT81), .A4(new_n415), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n413), .A2(KEYINPUT5), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n418), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G1gat), .B(G29gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT0), .ZN(new_n436));
  XNOR2_X1  g235(.A(G57gat), .B(G85gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT88), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n425), .B2(new_n433), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT6), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT6), .B1(new_n434), .B2(new_n439), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n433), .A3(new_n438), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT86), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(KEYINPUT86), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n265), .A2(new_n274), .ZN(new_n452));
  INV_X1    g251(.A(new_n256), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n281), .A2(new_n284), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n451), .B1(new_n454), .B2(new_n389), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT67), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT67), .B1(new_n262), .B2(new_n263), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n271), .A2(new_n272), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT27), .B(G183gat), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n459), .B(new_n259), .C1(new_n460), .C2(new_n258), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n458), .A2(new_n273), .B1(new_n461), .B2(new_n257), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n462), .A2(new_n256), .B1(new_n241), .B2(new_n250), .ZN(new_n463));
  INV_X1    g262(.A(new_n451), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n373), .B1(new_n455), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n468));
  OAI21_X1  g267(.A(new_n374), .B1(new_n251), .B2(new_n275), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n451), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT75), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n470), .B(new_n373), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT76), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT75), .B1(new_n454), .B2(new_n451), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n463), .A2(new_n472), .A3(new_n464), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n477), .A2(new_n478), .B1(new_n451), .B2(new_n469), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n479), .B2(new_n373), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n467), .B(new_n468), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G8gat), .B(G36gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G64gat), .B(G92gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n474), .A2(KEYINPUT76), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n476), .A3(new_n373), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n466), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT38), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n466), .B(new_n484), .C1(new_n486), .C2(new_n487), .ZN(new_n492));
  INV_X1    g291(.A(new_n484), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n488), .B2(new_n468), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n455), .A2(new_n373), .A3(new_n465), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n479), .B2(new_n373), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT38), .B1(new_n496), .B2(KEYINPUT37), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n449), .A2(new_n450), .A3(new_n491), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n412), .B1(new_n431), .B2(new_n418), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT39), .B1(new_n423), .B2(new_n413), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n438), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT39), .B(new_n412), .C1(new_n431), .C2(new_n418), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n504), .A2(KEYINPUT85), .A3(KEYINPUT40), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n467), .B(new_n493), .C1(new_n475), .C2(new_n480), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n467), .B1(new_n475), .B2(new_n480), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n484), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n487), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n467), .A4(new_n493), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT85), .B1(new_n504), .B2(KEYINPUT40), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n442), .B1(new_n504), .B2(KEYINPUT40), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n505), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n411), .B1(new_n499), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n398), .A2(new_n406), .A3(new_n400), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n406), .B1(new_n398), .B2(new_n400), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n518), .A2(new_n519), .A3(new_n409), .ZN(new_n520));
  INV_X1    g319(.A(new_n410), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g322(.A(new_n512), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n488), .A2(new_n493), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n512), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n434), .A2(new_n439), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n447), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n530), .A2(new_n440), .B1(new_n506), .B2(new_n507), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n319), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n508), .A2(new_n510), .A3(new_n535), .A4(new_n512), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n539), .A2(new_n450), .A3(new_n441), .A4(new_n444), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n311), .A2(new_n307), .A3(new_n313), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n408), .A2(new_n542), .A3(new_n410), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT89), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n408), .A2(new_n410), .A3(new_n309), .ZN(new_n545));
  OAI211_X1 g344(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n532), .C2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n536), .B1(new_n449), .B2(new_n450), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n408), .A2(new_n542), .A3(new_n410), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n425), .A2(new_n433), .A3(new_n438), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n552), .A2(new_n442), .A3(KEYINPUT6), .ZN(new_n553));
  INV_X1    g352(.A(new_n440), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n508), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT77), .B1(new_n510), .B2(new_n512), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n522), .A2(new_n557), .A3(new_n309), .A4(new_n527), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT90), .B1(new_n558), .B2(KEYINPUT35), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n534), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G183gat), .B(G211gat), .Z(new_n561));
  OR2_X1    g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G57gat), .A2(G64gat), .ZN(new_n563));
  AND2_X1   g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(KEYINPUT9), .ZN(new_n565));
  NOR2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n565), .A2(KEYINPUT98), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT98), .B1(new_n565), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n567), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT16), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(G1gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G15gat), .B(G22gat), .ZN(new_n586));
  MUX2_X1   g385(.A(G1gat), .B(new_n585), .S(new_n586), .Z(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(G8gat), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n573), .B2(new_n572), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT99), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n580), .A2(new_n581), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n583), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n592), .B1(new_n583), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n561), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  INV_X1    g397(.A(new_n561), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G134gat), .B(G162gat), .Z(new_n602));
  XOR2_X1   g401(.A(G43gat), .B(G50gat), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT15), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n606));
  OR3_X1    g405(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(G29gat), .A2(G36gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(KEYINPUT95), .A3(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n607), .B(KEYINPUT93), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n606), .B(KEYINPUT92), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n605), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT17), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT17), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n617), .A2(new_n624), .A3(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT7), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  AOI22_X1  g432(.A1(KEYINPUT8), .A2(new_n633), .B1(new_n627), .B2(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G99gat), .B(G106gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT101), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n635), .B(new_n637), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n626), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n635), .B(new_n637), .ZN(new_n640));
  AND2_X1   g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n622), .A2(new_n640), .B1(KEYINPUT41), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n639), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n645), .B2(new_n649), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n602), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  INV_X1    g453(.A(new_n602), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n572), .ZN(new_n659));
  INV_X1    g458(.A(new_n572), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n640), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n658), .B1(new_n662), .B2(KEYINPUT10), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n659), .A2(new_n661), .A3(KEYINPUT102), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n661), .A2(new_n664), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G230gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n292), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n662), .A2(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n673), .A2(new_n674), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n601), .A2(new_n657), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G113gat), .B(G141gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT11), .ZN(new_n685));
  INV_X1    g484(.A(G169gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n330), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n626), .A2(new_n589), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n622), .A2(new_n588), .ZN(new_n693));
  NAND2_X1  g492(.A1(G229gat), .A2(G233gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT96), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n693), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n626), .B2(new_n589), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(KEYINPUT96), .A3(new_n694), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT18), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(KEYINPUT18), .A3(new_n694), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n622), .B(new_n588), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n694), .B(KEYINPUT13), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n691), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n702), .A2(new_n690), .A3(new_n705), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n701), .B2(KEYINPUT97), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT18), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT96), .B1(new_n699), .B2(new_n694), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n588), .B1(new_n623), .B2(new_n625), .ZN(new_n713));
  INV_X1    g512(.A(new_n694), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n713), .A2(new_n698), .A3(new_n696), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT97), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n707), .B1(new_n710), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n560), .A2(new_n683), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n553), .A2(new_n554), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT103), .B(G1gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1324gat));
  INV_X1    g524(.A(new_n513), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT16), .B(G8gat), .Z(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT42), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(G8gat), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT42), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n732), .A2(KEYINPUT104), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT104), .B2(new_n732), .ZN(G1325gat));
  OAI21_X1  g535(.A(G15gat), .B1(new_n720), .B2(new_n319), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n314), .A2(G15gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n720), .B2(new_n738), .ZN(G1326gat));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n522), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT43), .B(G22gat), .Z(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1327gat));
  NAND2_X1  g541(.A1(new_n560), .A2(new_n657), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n682), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n601), .A2(new_n746), .A3(new_n719), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n657), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT35), .B1(new_n532), .B2(new_n545), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT90), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n752), .A2(new_n546), .A3(new_n544), .A4(new_n550), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n749), .B1(new_n753), .B2(new_n534), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n748), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n745), .A2(new_n755), .A3(KEYINPUT105), .A4(new_n748), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n722), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n748), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n762), .A2(G29gat), .A3(new_n722), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT45), .Z(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(G1328gat));
  OAI21_X1  g564(.A(G36gat), .B1(new_n760), .B2(new_n726), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n762), .A2(G36gat), .A3(new_n726), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1329gat));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  INV_X1    g569(.A(new_n319), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n758), .A2(new_n771), .A3(new_n759), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(G43gat), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n762), .A2(G43gat), .A3(new_n314), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n772), .B2(G43gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G43gat), .B1(new_n756), .B2(new_n319), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n775), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1330gat));
  OAI21_X1  g580(.A(G50gat), .B1(new_n756), .B2(new_n522), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n762), .A2(G50gat), .A3(new_n522), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(KEYINPUT48), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n758), .A2(new_n411), .A3(new_n759), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n786), .B2(G50gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G1331gat));
  INV_X1    g588(.A(new_n601), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n708), .B1(new_n716), .B2(new_n717), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n701), .A2(KEYINPUT97), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n716), .A2(new_n705), .A3(new_n702), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n691), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(new_n749), .A3(new_n682), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n753), .B2(new_n534), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n721), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g597(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT108), .ZN(new_n801));
  NOR2_X1   g600(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1333gat));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n771), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n314), .A2(G71gat), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n804), .A2(G71gat), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n796), .A2(new_n411), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g608(.A1(new_n601), .A2(new_n794), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n746), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n745), .A2(new_n755), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n745), .A2(new_n755), .A3(KEYINPUT109), .A4(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G85gat), .B1(new_n816), .B2(new_n722), .ZN(new_n817));
  INV_X1    g616(.A(new_n810), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n754), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n560), .A2(new_n657), .A3(new_n818), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n825), .A2(new_n627), .A3(new_n721), .A4(new_n682), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n817), .A2(new_n826), .ZN(G1336gat));
  OR2_X1    g626(.A1(new_n812), .A2(new_n726), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n628), .B1(new_n828), .B2(KEYINPUT112), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(KEYINPUT112), .B2(new_n828), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n746), .A2(G92gat), .A3(new_n726), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n814), .A2(new_n513), .A3(new_n815), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT51), .B1(new_n821), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n822), .A2(KEYINPUT111), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n821), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n835), .A2(G92gat), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n833), .B1(new_n834), .B2(new_n840), .ZN(G1337gat));
  OAI21_X1  g640(.A(G99gat), .B1(new_n816), .B2(new_n319), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n746), .A2(G99gat), .A3(new_n314), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT113), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n825), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(G1338gat));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n814), .A2(new_n411), .A3(new_n815), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G106gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n746), .A2(new_n522), .A3(G106gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n848), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G106gat), .B1(new_n812), .B2(new_n522), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n848), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n825), .A2(new_n851), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n825), .A2(KEYINPUT114), .A3(new_n851), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n847), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n854), .A2(new_n848), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n825), .A2(KEYINPUT114), .A3(new_n851), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT114), .B1(new_n825), .B2(new_n851), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n849), .A2(G106gat), .B1(new_n839), .B2(new_n851), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(KEYINPUT115), .C1(new_n848), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n867), .ZN(G1339gat));
  NOR4_X1   g667(.A1(new_n601), .A2(new_n719), .A3(new_n657), .A4(new_n682), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n669), .A2(new_n870), .A3(new_n672), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n667), .B1(new_n663), .B2(new_n665), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n671), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT54), .B1(new_n872), .B2(new_n671), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n678), .B(new_n871), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT55), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n673), .A2(KEYINPUT54), .A3(new_n873), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(KEYINPUT55), .A3(new_n678), .A4(new_n871), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n878), .A2(new_n880), .A3(new_n681), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n703), .A2(new_n704), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n714), .B1(new_n713), .B2(new_n698), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n688), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n791), .B2(new_n792), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n657), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n881), .A2(new_n719), .B1(new_n886), .B2(new_n682), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n657), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n869), .B1(new_n889), .B2(new_n601), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n722), .A2(new_n513), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n548), .ZN(new_n894));
  OAI21_X1  g693(.A(G113gat), .B1(new_n894), .B2(new_n794), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n890), .A2(new_n545), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n719), .A2(new_n210), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(G1340gat));
  NOR3_X1   g699(.A1(new_n894), .A2(new_n208), .A3(new_n746), .ZN(new_n901));
  AOI21_X1  g700(.A(G120gat), .B1(new_n896), .B2(new_n682), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n894), .B2(new_n601), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n220), .A3(new_n790), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1342gat));
  NOR3_X1   g705(.A1(new_n890), .A2(new_n749), .A3(new_n892), .ZN(new_n907));
  INV_X1    g706(.A(new_n545), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT68), .B(G134gat), .Z(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT56), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n222), .B1(new_n907), .B2(new_n548), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(G1343gat));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n771), .A2(new_n522), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n893), .A2(new_n344), .A3(new_n719), .A4(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n890), .B2(new_n522), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  INV_X1    g721(.A(new_n885), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n682), .B(new_n923), .C1(new_n710), .C2(new_n718), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n878), .A2(new_n880), .A3(new_n681), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n794), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n749), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n790), .B1(new_n927), .B2(new_n887), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n922), .B(new_n411), .C1(new_n928), .C2(new_n869), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n771), .A2(new_n892), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n921), .A2(new_n719), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT118), .ZN(new_n932));
  INV_X1    g731(.A(new_n930), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n411), .B1(new_n928), .B2(new_n869), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n920), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n719), .A4(new_n929), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n918), .B1(new_n938), .B2(G141gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n931), .A2(G141gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n917), .B1(new_n940), .B2(new_n916), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n914), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n941), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n344), .B1(new_n932), .B2(new_n937), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n943), .B(KEYINPUT119), .C1(new_n944), .C2(new_n918), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(G1344gat));
  AND2_X1   g745(.A1(new_n893), .A2(new_n915), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n345), .A3(new_n682), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G148gat), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n935), .A2(new_n929), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n682), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n934), .A2(KEYINPUT57), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n411), .B(new_n919), .C1(new_n928), .C2(new_n869), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n953), .A2(new_n682), .A3(new_n930), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n949), .B1(new_n955), .B2(G148gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n948), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(KEYINPUT120), .B(new_n948), .C1(new_n952), .C2(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1345gat));
  AOI21_X1  g760(.A(G155gat), .B1(new_n947), .B2(new_n790), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n790), .A2(G155gat), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT121), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n951), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT122), .ZN(G1346gat));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n350), .A3(new_n657), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n951), .A2(new_n657), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n350), .ZN(G1347gat));
  NOR3_X1   g768(.A1(new_n890), .A2(new_n721), .A3(new_n726), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n548), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n971), .A2(new_n686), .A3(new_n794), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n970), .A2(new_n908), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT123), .Z(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n719), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n972), .B1(new_n975), .B2(new_n686), .ZN(G1348gat));
  INV_X1    g775(.A(G176gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n977), .A3(new_n682), .ZN(new_n978));
  OAI21_X1  g777(.A(G176gat), .B1(new_n971), .B2(new_n746), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1349gat));
  NAND3_X1  g779(.A1(new_n973), .A2(new_n458), .A3(new_n790), .ZN(new_n981));
  OAI21_X1  g780(.A(G183gat), .B1(new_n971), .B2(new_n601), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g783(.A1(new_n974), .A2(new_n459), .A3(new_n657), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n548), .A3(new_n657), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(G190gat), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n987), .A2(new_n986), .A3(G190gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(G1351gat));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n915), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n330), .B1(new_n991), .B2(new_n794), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n319), .A2(new_n722), .A3(new_n513), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT124), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n794), .A2(new_n330), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n953), .A2(new_n954), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n992), .A2(new_n996), .ZN(G1352gat));
  NAND4_X1  g796(.A1(new_n970), .A2(new_n328), .A3(new_n682), .A4(new_n915), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  XOR2_X1   g798(.A(new_n999), .B(KEYINPUT125), .Z(new_n1000));
  NAND4_X1  g799(.A1(new_n953), .A2(new_n682), .A3(new_n954), .A4(new_n994), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G204gat), .ZN(new_n1002));
  OAI211_X1 g801(.A(new_n1000), .B(new_n1002), .C1(KEYINPUT62), .C2(new_n998), .ZN(G1353gat));
  INV_X1    g802(.A(new_n991), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1004), .A2(new_n334), .A3(new_n790), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n953), .A2(new_n790), .A3(new_n954), .A4(new_n994), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1006), .A2(G211gat), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(KEYINPUT63), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1005), .B1(new_n1010), .B2(new_n1011), .ZN(G1354gat));
  NAND3_X1  g811(.A1(new_n1004), .A2(new_n335), .A3(new_n657), .ZN(new_n1013));
  AND4_X1   g812(.A1(new_n657), .A2(new_n953), .A3(new_n954), .A4(new_n994), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n335), .B2(new_n1014), .ZN(G1355gat));
endmodule


