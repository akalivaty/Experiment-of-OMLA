//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n594, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n459), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT65), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT66), .ZN(G160));
  NOR2_X1   g048(.A1(new_n462), .A2(new_n463), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n459), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n459), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n477), .B2(G126), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n475), .A2(new_n488), .A3(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n475), .B2(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT72), .B1(new_n495), .B2(G543), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT71), .B(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n495), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n501));
  OAI211_X1 g076(.A(KEYINPUT72), .B(KEYINPUT5), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT69), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT69), .A2(G651), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT6), .A4(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT69), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT69), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n506), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n503), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT74), .B(G88), .Z(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n507), .A2(new_n508), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n514), .A2(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n521), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT75), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n525), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NOR3_X1   g110(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n503), .A2(new_n517), .A3(new_n514), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n517), .B1(new_n503), .B2(new_n514), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n539), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n503), .A2(G64), .ZN(new_n543));
  INV_X1    g118(.A(G77), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n499), .ZN(new_n545));
  INV_X1    g120(.A(new_n523), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(new_n546), .B1(G52), .B2(new_n534), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  AND2_X1   g124(.A1(new_n503), .A2(G56), .ZN(new_n550));
  AND2_X1   g125(.A1(G68), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n514), .A2(G43), .A3(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n539), .B2(G81), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI211_X1 g131(.A(KEYINPUT77), .B(new_n553), .C1(new_n539), .C2(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n565), .B1(new_n537), .B2(new_n538), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n516), .A2(KEYINPUT78), .A3(new_n518), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n566), .A2(new_n567), .A3(G91), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n503), .A2(KEYINPUT79), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n498), .A2(new_n576), .A3(new_n502), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n578), .B2(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n572), .B1(new_n579), .B2(new_n512), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT80), .B1(new_n568), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n498), .A2(new_n576), .A3(new_n502), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n576), .B1(new_n498), .B2(new_n502), .ZN(new_n583));
  OAI21_X1  g158(.A(G65), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n573), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n571), .B2(new_n570), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n566), .A2(new_n567), .A3(G91), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G299));
  AND2_X1   g166(.A1(new_n548), .A2(KEYINPUT81), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n548), .A2(KEYINPUT81), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G301));
  NAND2_X1  g170(.A1(new_n536), .A2(new_n540), .ZN(G286));
  NAND3_X1  g171(.A1(new_n566), .A2(new_n567), .A3(G87), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n503), .A2(G74), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n534), .B2(G49), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(G288));
  AOI22_X1  g175(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G48), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n601), .A2(new_n523), .B1(new_n602), .B2(new_n525), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n566), .A2(new_n567), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G86), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n523), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT83), .B(G47), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n608), .A2(new_n609), .B1(new_n534), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT84), .B(G85), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n539), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n611), .B(new_n613), .C1(new_n609), .C2(new_n608), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT85), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n575), .B2(new_n577), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n617), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(G66), .B1(new_n582), .B2(new_n583), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n623), .A2(KEYINPUT86), .A3(new_n620), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n622), .A2(G651), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n534), .A2(G54), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n566), .A2(new_n567), .A3(G92), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT10), .A4(G92), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n616), .B1(G868), .B2(new_n632), .ZN(G284));
  OAI21_X1  g208(.A(new_n616), .B1(G868), .B2(new_n632), .ZN(G321));
  NAND2_X1  g209(.A1(G286), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n590), .B2(G868), .ZN(G297));
  OAI21_X1  g211(.A(new_n635), .B1(new_n590), .B2(G868), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n632), .B1(new_n638), .B2(G860), .ZN(G148));
  INV_X1    g214(.A(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n558), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n630), .A2(new_n631), .ZN(new_n642));
  INV_X1    g217(.A(new_n626), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n624), .A2(G651), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n622), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n646), .A2(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n641), .B1(new_n647), .B2(new_n640), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n464), .A2(new_n460), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT12), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  AOI22_X1  g229(.A1(G123), .A2(new_n477), .B1(new_n475), .B2(G135), .ZN(new_n655));
  OAI21_X1  g230(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n656));
  INV_X1    g231(.A(G111), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n656), .A2(KEYINPUT88), .B1(new_n657), .B2(G2105), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(KEYINPUT88), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2096), .Z(new_n661));
  OAI211_X1 g236(.A(new_n654), .B(new_n661), .C1(G2100), .C2(new_n652), .ZN(G156));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT89), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(KEYINPUT14), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT16), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  NOR2_X1   g257(.A1(G2072), .A2(G2078), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n442), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(KEYINPUT17), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n680), .B(new_n681), .C1(new_n442), .C2(new_n683), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT18), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2096), .B(G2100), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1956), .B(G2474), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT20), .ZN(new_n702));
  INV_X1    g277(.A(new_n700), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n705), .B(new_n704), .S(new_n697), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(G229));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G5), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G171), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G1961), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n716), .A2(G21), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G286), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1966), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G160), .A2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n725), .B2(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT101), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n723), .B(new_n731), .C1(new_n722), .C2(new_n721), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G33), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT99), .B(KEYINPUT25), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(new_n459), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n737), .B(new_n739), .C1(G139), .C2(new_n475), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n733), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT30), .B(G28), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n743), .A2(new_n733), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n742), .B(new_n746), .C1(new_n733), .C2(new_n660), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n741), .A2(G2072), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n733), .A2(G32), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n477), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n460), .A2(G105), .ZN(new_n754));
  INV_X1    g329(.A(G141), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n465), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(new_n733), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n733), .A2(G26), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT28), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n475), .A2(G140), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n477), .A2(G128), .ZN(new_n765));
  OR2_X1    g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n747), .A2(new_n748), .A3(new_n761), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G27), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n773), .A2(KEYINPUT102), .A3(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT102), .B1(new_n773), .B2(G29), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G164), .C2(new_n733), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G2078), .Z(new_n777));
  OAI211_X1 g352(.A(new_n772), .B(new_n777), .C1(new_n729), .C2(new_n728), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n733), .A2(G35), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT103), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n482), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT29), .ZN(new_n782));
  INV_X1    g357(.A(G2090), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n782), .A2(new_n783), .B1(G1961), .B2(new_n718), .ZN(new_n784));
  AOI21_X1  g359(.A(KEYINPUT104), .B1(new_n782), .B2(new_n783), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n782), .A2(KEYINPUT104), .A3(new_n783), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n778), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n646), .A2(G16), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G4), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1348), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G1348), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n732), .A2(new_n787), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G19), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n559), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1341), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n716), .A2(G20), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT23), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n590), .B2(new_n716), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1956), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n794), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n597), .A2(new_n599), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n808));
  NAND2_X1  g383(.A1(G288), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G23), .B(new_n810), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT33), .B(G1976), .Z(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n605), .A2(new_n716), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G6), .B2(new_n716), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n716), .A2(G22), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G166), .B2(new_n716), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1971), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n818), .A2(new_n820), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n733), .A2(G25), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n829));
  INV_X1    g404(.A(G107), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(G2105), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT94), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G119), .B2(new_n477), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n475), .A2(G131), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT93), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT95), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n828), .B1(new_n841), .B2(new_n733), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G1986), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n716), .A2(G24), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G290), .B2(G16), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n844), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n845), .B2(new_n847), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n827), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n814), .A2(new_n816), .A3(new_n826), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT34), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n805), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n805), .A3(new_n852), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n804), .B1(new_n854), .B2(new_n855), .ZN(G311));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n803), .B1(new_n857), .B2(new_n853), .ZN(G150));
  NOR2_X1   g433(.A1(new_n646), .A2(new_n638), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n539), .A2(G93), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n862), .A2(new_n523), .B1(new_n863), .B2(new_n525), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n559), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n558), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n860), .B(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n865), .A2(new_n872), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  XNOR2_X1  g452(.A(new_n840), .B(KEYINPUT105), .ZN(new_n878));
  INV_X1    g453(.A(new_n651), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n475), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n477), .A2(G130), .ZN(new_n884));
  OR2_X1    g459(.A1(G106), .A2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n885), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n880), .A2(new_n889), .A3(new_n881), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n491), .B(new_n768), .ZN(new_n893));
  INV_X1    g468(.A(new_n757), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n740), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G160), .B(new_n660), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n901));
  INV_X1    g476(.A(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n891), .B2(new_n896), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n888), .A2(new_n902), .A3(new_n890), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g484(.A1(new_n810), .A2(new_n605), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n807), .A2(G305), .A3(new_n809), .ZN(new_n911));
  XNOR2_X1  g486(.A(G290), .B(G303), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT42), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(new_n911), .ZN(new_n919));
  INV_X1    g494(.A(new_n912), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT109), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n916), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n918), .A2(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT110), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n869), .A2(new_n647), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n869), .A2(new_n647), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n581), .A2(KEYINPUT107), .A3(new_n589), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n632), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n646), .A2(KEYINPUT107), .A3(new_n581), .A4(new_n589), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n930), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n936), .B2(new_n937), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT108), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n929), .A2(new_n930), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n926), .A2(new_n928), .A3(new_n939), .A4(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n926), .A2(new_n928), .B1(new_n939), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(G868), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n865), .A2(G868), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(G295));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n952), .A2(new_n956), .A3(new_n954), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n926), .A2(new_n928), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n948), .A2(new_n939), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n640), .B1(new_n960), .B2(new_n949), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT111), .B1(new_n961), .B2(new_n953), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n962), .ZN(G331));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g539(.A(G168), .B1(new_n592), .B2(new_n593), .ZN(new_n965));
  NAND2_X1  g540(.A1(G286), .A2(new_n548), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n868), .A3(new_n866), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n558), .A2(new_n867), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n558), .A2(new_n867), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n965), .B(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n938), .A2(KEYINPUT41), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n946), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n947), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n937), .A3(new_n936), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n980), .B2(new_n927), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n972), .A2(new_n938), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n943), .A2(new_n947), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n972), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n918), .A2(new_n923), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT43), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n941), .A2(new_n942), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n979), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  AOI21_X1  g564(.A(G37), .B1(new_n989), .B2(new_n927), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n977), .A2(new_n985), .A3(new_n979), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n964), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n978), .B1(new_n943), .B2(new_n947), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n927), .B1(new_n995), .B2(new_n982), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n991), .A3(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n998), .A2(KEYINPUT43), .B1(new_n986), .B2(new_n990), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n964), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n491), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n472), .A2(G40), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1003), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(KEYINPUT126), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT126), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1005), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n768), .B(new_n770), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n894), .B(new_n1014), .C1(KEYINPUT46), .C2(new_n1006), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1010), .A2(new_n1011), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT47), .Z(new_n1017));
  NAND3_X1  g592(.A1(new_n1005), .A2(G1996), .A3(new_n894), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT112), .Z(new_n1019));
  AOI21_X1  g594(.A(new_n1014), .B1(new_n1006), .B2(new_n757), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n841), .A2(new_n843), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT125), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1021), .A2(new_n1023), .B1(G2067), .B2(new_n768), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(new_n1005), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n840), .B(new_n843), .Z(new_n1026));
  AOI21_X1  g601(.A(new_n1021), .B1(new_n1005), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1012), .A2(G290), .A3(G1986), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT48), .Z(new_n1029));
  AOI211_X1 g604(.A(new_n1017), .B(new_n1025), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n472), .A2(G40), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1003), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n605), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT115), .B(G86), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n519), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(G1981), .B1(new_n1037), .B2(new_n603), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1033), .B1(new_n1041), .B2(KEYINPUT49), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(KEYINPUT49), .B2(new_n1041), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n806), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1035), .B(KEYINPUT117), .Z(new_n1046));
  AOI21_X1  g621(.A(new_n1033), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n810), .A2(new_n1044), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n1048), .B2(new_n1033), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1033), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1044), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1043), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1031), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1001), .B1(new_n492), .B2(new_n493), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(KEYINPUT50), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n783), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(KEYINPUT113), .A3(new_n1061), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1002), .A2(new_n1061), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n1004), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1971), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1060), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1055), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT114), .B1(new_n1073), .B2(new_n1060), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G303), .A2(G8), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1075), .B(KEYINPUT55), .Z(new_n1076));
  AND3_X1   g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1047), .B1(new_n1054), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1004), .B1(new_n1002), .B2(new_n1061), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n722), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1058), .A2(new_n729), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1055), .B1(new_n1084), .B2(G168), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(G286), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1068), .B2(G2078), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1058), .A2(G1961), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G2078), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1080), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n594), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1087), .A2(new_n1089), .B1(KEYINPUT62), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n568), .A2(new_n580), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT57), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1004), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1057), .B2(KEYINPUT50), .ZN(new_n1103));
  INV_X1    g678(.A(G1956), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1101), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1058), .A2(G1348), .B1(G2067), .B2(new_n1032), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1110), .A2(new_n632), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(new_n632), .ZN(new_n1116));
  OR3_X1    g691(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1116), .A2(new_n1117), .B1(new_n1114), .B2(new_n1110), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT58), .B(G1341), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1032), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT121), .Z(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(G1996), .B2(new_n1068), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n559), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1108), .A2(KEYINPUT61), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(KEYINPUT59), .A3(new_n559), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1108), .A2(KEYINPUT61), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1112), .B1(new_n1118), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1066), .A2(new_n1095), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1092), .A2(KEYINPUT124), .B1(new_n1079), .B2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1091), .B(new_n1133), .C1(KEYINPUT124), .C2(new_n1092), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1098), .B(new_n1131), .C1(new_n594), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1097), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1136), .A2(G301), .B1(new_n1134), .B2(G171), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1137), .B2(new_n1131), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1099), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1103), .A2(G2090), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1073), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1076), .B1(new_n1141), .B2(G8), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1077), .A2(new_n1053), .A3(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1097), .A2(KEYINPUT62), .A3(new_n594), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1078), .B1(new_n1139), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1148));
  NOR3_X1   g723(.A1(new_n1084), .A2(new_n1055), .A3(G286), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(KEYINPUT63), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1077), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1076), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1053), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1053), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1152), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1150), .B1(new_n1158), .B2(KEYINPUT120), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n1152), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1147), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G290), .B(new_n845), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1027), .B1(new_n1012), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1030), .B1(new_n1162), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g740(.A(G319), .B(new_n693), .C1(new_n677), .C2(new_n678), .ZN(new_n1167));
  INV_X1    g741(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n714), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n900), .B1(new_n892), .B2(new_n896), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n896), .B2(new_n892), .ZN(new_n1172));
  INV_X1    g746(.A(new_n907), .ZN(new_n1173));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n999), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1169), .B1(new_n904), .B2(new_n907), .ZN(new_n1177));
  INV_X1    g751(.A(KEYINPUT43), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n981), .B2(new_n991), .ZN(new_n1179));
  AND3_X1   g753(.A1(new_n990), .A2(new_n991), .A3(new_n1178), .ZN(new_n1180));
  OAI211_X1 g754(.A(new_n1176), .B(new_n1177), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AND2_X1   g755(.A1(new_n1175), .A2(new_n1181), .ZN(G308));
  NAND2_X1  g756(.A1(new_n1175), .A2(new_n1181), .ZN(G225));
endmodule


