//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944;
  XNOR2_X1  g000(.A(KEYINPUT24), .B(G110), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G119), .B(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n191), .B2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT73), .B1(new_n193), .B2(G128), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI22_X1  g010(.A1(new_n189), .A2(new_n190), .B1(new_n196), .B2(G110), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n200), .A2(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n203), .B1(new_n206), .B2(new_n199), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT74), .A3(new_n202), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT74), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n201), .A2(new_n209), .A3(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(G110), .B2(new_n196), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n189), .A2(new_n190), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n205), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT22), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(G137), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n217), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G217), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G234), .B2(new_n223), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n222), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n231), .B2(new_n226), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT32), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT11), .A2(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT11), .A2(G134), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(G137), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT64), .B(G137), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n239), .B(new_n240), .C1(new_n238), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT11), .A3(G134), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(KEYINPUT65), .A3(new_n240), .A4(new_n239), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT66), .B1(new_n249), .B2(G134), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n241), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(G134), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n252), .A2(KEYINPUT67), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT67), .B1(new_n252), .B2(new_n259), .ZN(new_n261));
  XNOR2_X1  g075(.A(G143), .B(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G128), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n191), .A2(new_n203), .A3(G143), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(G146), .C1(new_n191), .C2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n260), .A2(new_n261), .A3(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n250), .A2(new_n239), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n252), .B1(new_n240), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(KEYINPUT0), .B(G128), .Z(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n262), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n236), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n193), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G119), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT2), .B(G113), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n252), .A2(new_n259), .A3(new_n268), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT68), .B(new_n236), .C1(new_n270), .C2(new_n278), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n281), .A2(new_n287), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n288), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(G101), .ZN(new_n295));
  NOR2_X1   g109(.A1(G237), .A2(G953), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G210), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n295), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n235), .B1(new_n301), .B2(KEYINPUT31), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT69), .B(new_n303), .C1(new_n291), .C2(new_n300), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n291), .A2(new_n303), .A3(new_n300), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n293), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n292), .A2(KEYINPUT28), .A3(new_n287), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n287), .ZN(new_n310));
  INV_X1    g124(.A(new_n270), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n277), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n299), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n305), .A2(new_n313), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n302), .A2(new_n304), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G472), .A2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n234), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n301), .A2(KEYINPUT31), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT69), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n305), .A2(new_n313), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n301), .A2(new_n235), .A3(KEYINPUT31), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT32), .A3(new_n316), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n316), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT70), .A3(new_n234), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT71), .ZN(new_n330));
  INV_X1    g144(.A(new_n293), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n291), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n299), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n309), .A2(new_n312), .A3(new_n299), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n292), .A2(new_n287), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n309), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n299), .A2(new_n334), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n330), .B1(new_n342), .B2(G472), .ZN(new_n343));
  INV_X1    g157(.A(G472), .ZN(new_n344));
  AOI211_X1 g158(.A(KEYINPUT71), .B(new_n344), .C1(new_n336), .C2(new_n341), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n233), .B1(new_n329), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G104), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n350), .B(new_n353), .C1(G104), .C2(new_n352), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(G101), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(G101), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n358), .A3(G101), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n287), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n352), .A2(G104), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n349), .A2(G107), .ZN(new_n364));
  OAI21_X1  g178(.A(G101), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n285), .A2(new_n286), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT5), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G113), .B1(new_n282), .B2(KEYINPUT5), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n357), .A2(KEYINPUT81), .A3(new_n287), .A4(new_n359), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT82), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT83), .B1(new_n377), .B2(KEYINPUT6), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n374), .A2(new_n379), .A3(new_n380), .A4(new_n376), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n276), .A2(G125), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n269), .B2(G125), .ZN(new_n384));
  INV_X1    g198(.A(G224), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G953), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n384), .B(new_n386), .Z(new_n387));
  OR2_X1    g201(.A1(new_n374), .A2(new_n376), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n382), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n376), .B(KEYINPUT84), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n391), .B(KEYINPUT8), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n366), .A2(new_n371), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n368), .B(KEYINPUT85), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n367), .B1(new_n394), .B2(new_n370), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n366), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n387), .B1(KEYINPUT7), .B2(new_n386), .ZN(new_n398));
  OR3_X1    g212(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n386), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n388), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n223), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G210), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n348), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(KEYINPUT86), .A3(new_n403), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n348), .B1(new_n403), .B2(KEYINPUT86), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n390), .A2(new_n223), .A3(new_n400), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G221), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT9), .B(G234), .Z(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n223), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G469), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n366), .A2(new_n269), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n355), .A2(new_n268), .A3(new_n365), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n419), .A2(KEYINPUT79), .A3(KEYINPUT12), .A4(new_n272), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n419), .A2(new_n272), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(KEYINPUT12), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n357), .A2(new_n276), .A3(new_n359), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n276), .A4(new_n359), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n430));
  AOI22_X1  g244(.A1(new_n428), .A2(new_n429), .B1(new_n418), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n272), .ZN(new_n432));
  INV_X1    g246(.A(new_n418), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(KEYINPUT10), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n218), .A2(G227), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n438), .B(new_n439), .Z(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT76), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n432), .B1(new_n431), .B2(new_n435), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n436), .A3(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n416), .B1(new_n446), .B2(new_n223), .ZN(new_n447));
  INV_X1    g261(.A(new_n440), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n425), .A2(new_n436), .A3(new_n440), .ZN(new_n451));
  AOI211_X1 g265(.A(G469), .B(G902), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n415), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n451), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n416), .A3(new_n223), .ZN(new_n456));
  NAND2_X1  g270(.A1(G469), .A2(G902), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n456), .B(new_n457), .C1(new_n416), .C2(new_n446), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n415), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n296), .A2(G143), .A3(G214), .ZN(new_n462));
  AOI21_X1  g276(.A(G143), .B1(new_n296), .B2(G214), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n240), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT89), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n467), .A2(new_n466), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n471), .A3(new_n466), .A4(new_n467), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n211), .A2(new_n469), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT18), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n464), .B1(new_n474), .B2(new_n240), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n200), .B(new_n203), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(new_n476), .C1(new_n467), .C2(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G113), .B(G122), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(new_n349), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT90), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n473), .A2(new_n483), .A3(new_n480), .A4(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n223), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G475), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n200), .B(KEYINPUT19), .Z(new_n490));
  OAI21_X1  g304(.A(new_n202), .B1(new_n490), .B2(G146), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n465), .A2(new_n467), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n477), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n481), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n482), .A2(new_n484), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR4_X1   g311(.A1(new_n497), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G475), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n223), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT20), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n498), .B1(new_n503), .B2(KEYINPUT91), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT20), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n489), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G128), .B(G143), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n255), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n283), .A2(KEYINPUT14), .A3(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(G116), .B(G122), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(G107), .B(new_n510), .C1(new_n512), .C2(KEYINPUT14), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n509), .B(new_n513), .C1(G107), .C2(new_n512), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(KEYINPUT13), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n266), .A2(G128), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(G134), .C1(KEYINPUT13), .C2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n511), .B(new_n352), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(new_n255), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n413), .A2(G217), .A3(new_n218), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n521), .B(new_n522), .Z(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(G902), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT92), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n524), .B(KEYINPUT92), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n507), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT93), .B(G952), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n535), .A2(G902), .A3(G953), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n411), .A2(new_n461), .A3(new_n532), .A4(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n347), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(G101), .ZN(G3));
  NAND2_X1  g359(.A1(new_n324), .A2(new_n223), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G472), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n232), .A2(new_n461), .A3(new_n547), .A4(new_n327), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OR3_X1    g363(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n403), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n401), .A2(new_n403), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n401), .A2(KEYINPUT95), .A3(new_n403), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT94), .B1(new_n401), .B2(new_n403), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n550), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n409), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n526), .A2(new_n223), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n524), .A2(new_n526), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT33), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n521), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n523), .B(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n558), .B(new_n560), .C1(new_n564), .C2(G478), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n507), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n557), .A2(new_n540), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n549), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT34), .B(G104), .Z(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G6));
  INV_X1    g384(.A(new_n557), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n489), .B(KEYINPUT97), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  AOI21_X1  g387(.A(G475), .B1(new_n485), .B2(new_n499), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n223), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n498), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n572), .A2(new_n530), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n540), .B(KEYINPUT98), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n549), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G107), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G9));
  NAND2_X1  g396(.A1(new_n231), .A2(new_n226), .ZN(new_n583));
  INV_X1    g397(.A(new_n221), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n217), .B(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n223), .C1(new_n225), .C2(G234), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n547), .A2(new_n327), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n542), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT37), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G110), .ZN(G12));
  NAND2_X1  g406(.A1(new_n329), .A2(new_n346), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n588), .A2(new_n557), .ZN(new_n594));
  INV_X1    g408(.A(G900), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n537), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n536), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n577), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n593), .A2(new_n594), .A3(new_n461), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G128), .ZN(G30));
  OAI21_X1  g415(.A(new_n299), .B1(new_n338), .B2(new_n293), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT99), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n301), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n344), .B1(new_n604), .B2(new_n223), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n329), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n489), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n503), .A2(new_n498), .A3(KEYINPUT91), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n574), .A2(new_n573), .A3(new_n223), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n575), .B2(new_n505), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n530), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n408), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT38), .A4(new_n407), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n613), .A2(new_n615), .A3(new_n409), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n607), .A2(new_n588), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT100), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n597), .B(KEYINPUT39), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n461), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT101), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n461), .A2(new_n625), .A3(new_n622), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(KEYINPUT40), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n461), .B2(new_n622), .ZN(new_n629));
  AOI211_X1 g443(.A(KEYINPUT101), .B(new_n621), .C1(new_n454), .C2(new_n460), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n583), .A2(new_n587), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n329), .B2(new_n606), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n618), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n620), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  INV_X1    g453(.A(new_n565), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n612), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n598), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n593), .A2(new_n594), .A3(new_n461), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G146), .ZN(G48));
  AOI21_X1  g459(.A(new_n416), .B1(new_n455), .B2(new_n223), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n452), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n415), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT102), .Z(new_n649));
  NAND3_X1  g463(.A1(new_n347), .A2(new_n567), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT41), .B(G113), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  NAND3_X1  g466(.A1(new_n347), .A2(new_n579), .A3(new_n649), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G116), .ZN(G18));
  NOR4_X1   g468(.A1(new_n507), .A2(new_n648), .A3(new_n540), .A4(new_n531), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n593), .A2(new_n594), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G119), .ZN(G21));
  OAI211_X1 g471(.A(new_n320), .B(new_n305), .C1(new_n298), .C2(new_n339), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n316), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT103), .B1(new_n546), .B2(G472), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n661), .B(new_n344), .C1(new_n324), .C2(new_n223), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n232), .B(new_n659), .C1(new_n660), .C2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n571), .A2(new_n578), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n613), .A4(new_n649), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT104), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(G122), .Z(G24));
  OAI21_X1  g482(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n588), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n642), .A2(new_n557), .A3(new_n648), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G125), .ZN(G27));
  XNOR2_X1  g487(.A(new_n458), .B(KEYINPUT105), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n643), .A2(new_n415), .A3(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n318), .B(new_n325), .C1(new_n343), .C2(new_n345), .ZN(new_n676));
  INV_X1    g490(.A(new_n409), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n408), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n232), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n674), .A2(new_n415), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n642), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n347), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n240), .ZN(G33));
  NOR2_X1   g500(.A1(new_n681), .A2(new_n597), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n347), .A2(new_n577), .A3(new_n678), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G134), .ZN(G36));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n507), .B2(new_n640), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n612), .A2(KEYINPUT43), .A3(new_n565), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n589), .A3(new_n634), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n449), .A2(new_n443), .A3(new_n448), .ZN(new_n698));
  INV_X1    g512(.A(new_n441), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n425), .B2(new_n436), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n442), .A2(KEYINPUT45), .A3(new_n445), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n702), .A3(G469), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n457), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT106), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n703), .A2(KEYINPUT46), .A3(new_n457), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n704), .A2(new_n709), .A3(new_n705), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n456), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n415), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n621), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n693), .A2(new_n589), .A3(new_n634), .A4(KEYINPUT44), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n678), .B(KEYINPUT107), .Z(new_n715));
  NAND4_X1  g529(.A1(new_n696), .A2(new_n713), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G137), .ZN(G39));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n711), .A2(KEYINPUT47), .A3(new_n415), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n642), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n593), .A2(new_n232), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n678), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G140), .ZN(G42));
  INV_X1    g538(.A(new_n461), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n329), .B2(new_n346), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n572), .A2(new_n531), .A3(new_n576), .A4(new_n597), .ZN(new_n727));
  INV_X1    g541(.A(new_n669), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n726), .A2(new_n727), .B1(new_n728), .B2(new_n682), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n634), .A2(new_n678), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n688), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(new_n688), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n683), .A2(new_n684), .ZN(new_n736));
  INV_X1    g550(.A(new_n680), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n593), .A2(new_n232), .A3(new_n543), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n566), .A2(KEYINPUT109), .B1(new_n531), .B2(new_n612), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n612), .A2(KEYINPUT109), .A3(new_n531), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n411), .B(new_n578), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n548), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n739), .A2(new_n744), .A3(new_n590), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n653), .A2(new_n666), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n650), .A2(new_n656), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n738), .A2(new_n745), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n726), .B(new_n594), .C1(new_n599), .C2(new_n643), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n557), .A2(new_n530), .A3(new_n612), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n635), .A2(new_n687), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n735), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n672), .A3(new_n751), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n752), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT53), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n758), .A2(new_n735), .A3(new_n761), .A4(new_n748), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT54), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n764));
  INV_X1    g578(.A(new_n678), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n765), .B2(new_n648), .ZN(new_n766));
  INV_X1    g580(.A(new_n536), .ZN(new_n767));
  INV_X1    g581(.A(new_n648), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n678), .A2(KEYINPUT115), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n607), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n232), .A3(new_n641), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n534), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n693), .A2(new_n767), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n663), .A2(new_n774), .A3(new_n648), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n773), .B1(new_n571), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n647), .B(KEYINPUT112), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n719), .B(new_n720), .C1(new_n415), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n663), .A2(new_n774), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n715), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT113), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n615), .A2(new_n616), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n409), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n775), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n782), .B1(new_n775), .B2(new_n785), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT51), .B(new_n780), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n770), .B1(new_n691), .B2(new_n692), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n670), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n771), .A2(new_n232), .A3(new_n612), .A4(new_n640), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n776), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n793), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n787), .A2(KEYINPUT114), .A3(new_n788), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n775), .A2(new_n785), .ZN(new_n798));
  INV_X1    g612(.A(new_n782), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n797), .B1(new_n800), .B2(new_n786), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n795), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n795), .B(KEYINPUT116), .C1(new_n796), .C2(new_n801), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n780), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n794), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n761), .B1(new_n754), .B2(new_n759), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n758), .A2(new_n735), .A3(new_n748), .A4(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n763), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n676), .A2(new_n232), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n790), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT48), .Z(new_n816));
  OAI22_X1  g630(.A1(new_n813), .A2(new_n816), .B1(G952), .B2(G953), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n507), .A2(new_n677), .A3(new_n640), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n232), .A3(new_n415), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n784), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n605), .B1(new_n326), .B2(new_n328), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n647), .B(KEYINPUT49), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(G75));
  NAND4_X1  g640(.A1(new_n650), .A2(new_n653), .A3(new_n666), .A4(new_n656), .ZN(new_n827));
  INV_X1    g641(.A(new_n590), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n544), .B(new_n828), .C1(new_n548), .C2(new_n743), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n827), .A2(new_n685), .A3(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n600), .A2(new_n644), .A3(new_n672), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT52), .A4(new_n751), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n833), .A3(new_n734), .A4(new_n732), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n757), .A2(new_n752), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n832), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n735), .A2(new_n748), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n761), .A3(new_n835), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n839), .A3(G210), .A4(G902), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n382), .A2(new_n389), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(new_n387), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT55), .Z(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n840), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n840), .B2(new_n841), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n218), .A2(G952), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G51));
  XOR2_X1   g663(.A(new_n457), .B(KEYINPUT57), .Z(new_n850));
  AND3_X1   g664(.A1(new_n837), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT54), .B1(new_n837), .B2(new_n839), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n455), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n837), .A2(G902), .A3(new_n839), .ZN(new_n855));
  INV_X1    g669(.A(new_n703), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n848), .B1(new_n854), .B2(new_n857), .ZN(G54));
  NAND3_X1  g672(.A1(new_n855), .A2(KEYINPUT58), .A3(G475), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n497), .ZN(new_n860));
  INV_X1    g674(.A(new_n848), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(KEYINPUT58), .A3(G475), .A4(new_n500), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G60));
  INV_X1    g677(.A(new_n564), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n558), .B(KEYINPUT59), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n866), .C1(new_n851), .C2(new_n852), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n763), .B2(new_n812), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n861), .B(new_n867), .C1(new_n868), .C2(new_n864), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(G63));
  XNOR2_X1  g684(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n225), .A2(new_n223), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n837), .A2(new_n839), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n222), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n586), .B(KEYINPUT120), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n837), .A2(new_n839), .A3(new_n875), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n861), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(KEYINPUT61), .A3(new_n861), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(G66));
  OAI21_X1  g699(.A(G953), .B1(new_n538), .B2(new_n385), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n827), .A2(new_n829), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n842), .B1(G898), .B2(new_n218), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(G69));
  AOI21_X1  g704(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n281), .A2(new_n289), .A3(new_n290), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(new_n490), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(G900), .A2(G953), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n713), .A2(new_n814), .A3(new_n750), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT124), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n723), .A2(new_n716), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n749), .A2(new_n672), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n685), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n896), .A2(KEYINPUT124), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n900), .A3(new_n688), .A4(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n894), .B(new_n895), .C1(new_n902), .C2(G953), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n891), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n636), .B1(new_n635), .B2(new_n618), .ZN(new_n907));
  NOR4_X1   g721(.A1(new_n823), .A2(KEYINPUT100), .A3(new_n634), .A4(new_n617), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n632), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT62), .B1(new_n909), .B2(new_n899), .ZN(new_n910));
  INV_X1    g724(.A(new_n740), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n623), .B1(new_n911), .B2(new_n741), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n347), .A3(new_n678), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n723), .A2(new_n716), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n638), .A2(new_n831), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n910), .A2(KEYINPUT121), .A3(new_n916), .A4(new_n914), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n218), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n893), .ZN(new_n924));
  AOI21_X1  g738(.A(G953), .B1(new_n919), .B2(new_n920), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT122), .B1(new_n925), .B2(new_n894), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n906), .B1(new_n927), .B2(new_n903), .ZN(new_n928));
  INV_X1    g742(.A(new_n903), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n929), .B(new_n905), .C1(new_n924), .C2(new_n926), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G72));
  XNOR2_X1  g745(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n344), .A2(new_n223), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n932), .B(new_n933), .Z(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n333), .B2(new_n301), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT127), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n760), .B2(new_n762), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n332), .B(KEYINPUT126), .Z(new_n938));
  NOR3_X1   g752(.A1(new_n902), .A2(new_n827), .A3(new_n829), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n299), .B(new_n938), .C1(new_n939), .C2(new_n934), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n861), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n919), .A2(new_n887), .A3(new_n920), .ZN(new_n942));
  INV_X1    g756(.A(new_n934), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n298), .B2(new_n944), .ZN(G57));
endmodule


