

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721;

  XNOR2_X1 U370 ( .A(n437), .B(G134), .ZN(n458) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n487) );
  INV_X1 U372 ( .A(G146), .ZN(n439) );
  NOR2_X1 U373 ( .A1(G902), .A2(n600), .ZN(n498) );
  NOR2_X2 U374 ( .A1(n716), .A2(n393), .ZN(n374) );
  NOR2_X2 U375 ( .A1(n645), .A2(n565), .ZN(n566) );
  NOR2_X2 U376 ( .A1(n662), .A2(n661), .ZN(n509) );
  XNOR2_X2 U377 ( .A(n549), .B(n548), .ZN(n557) );
  NOR2_X2 U378 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X2 U379 ( .A(n511), .B(KEYINPUT1), .ZN(n555) );
  NOR2_X2 U380 ( .A1(n526), .A2(n522), .ZN(n621) );
  XOR2_X2 U381 ( .A(KEYINPUT6), .B(n568), .Z(n554) );
  NOR2_X1 U382 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U383 ( .A1(n556), .A2(n646), .ZN(n569) );
  XNOR2_X1 U384 ( .A(n471), .B(n363), .ZN(n643) );
  XNOR2_X1 U385 ( .A(n704), .B(n439), .ZN(n496) );
  XNOR2_X1 U386 ( .A(n409), .B(n455), .ZN(n697) );
  XNOR2_X1 U387 ( .A(n396), .B(KEYINPUT81), .ZN(n395) );
  INV_X2 U388 ( .A(G128), .ZN(n401) );
  XOR2_X1 U389 ( .A(KEYINPUT67), .B(G101), .Z(n491) );
  AND2_X2 U390 ( .A1(n585), .A2(n584), .ZN(n349) );
  XOR2_X2 U391 ( .A(n532), .B(KEYINPUT38), .Z(n659) );
  BUF_X2 U392 ( .A(n518), .Z(n532) );
  NAND2_X1 U393 ( .A1(n383), .A2(n382), .ZN(n381) );
  AND2_X1 U394 ( .A1(n533), .A2(n618), .ZN(n383) );
  NOR2_X1 U395 ( .A1(n619), .A2(n524), .ZN(n525) );
  NOR2_X1 U396 ( .A1(n643), .A2(n642), .ZN(n646) );
  XNOR2_X1 U397 ( .A(n381), .B(n380), .ZN(n405) );
  XNOR2_X1 U398 ( .A(n439), .B(G125), .ZN(n442) );
  XNOR2_X1 U399 ( .A(n430), .B(KEYINPUT93), .ZN(n413) );
  XNOR2_X1 U400 ( .A(n391), .B(n351), .ZN(n527) );
  OR2_X1 U401 ( .A1(n592), .A2(G902), .ZN(n391) );
  XNOR2_X1 U402 ( .A(n441), .B(n398), .ZN(n397) );
  OR2_X1 U403 ( .A1(n681), .A2(G902), .ZN(n399) );
  INV_X1 U404 ( .A(G472), .ZN(n497) );
  XNOR2_X1 U405 ( .A(G110), .B(G104), .ZN(n415) );
  XNOR2_X1 U406 ( .A(n442), .B(n390), .ZN(n703) );
  XNOR2_X1 U407 ( .A(G140), .B(KEYINPUT10), .ZN(n390) );
  XNOR2_X1 U408 ( .A(n407), .B(n515), .ZN(n541) );
  NOR2_X1 U409 ( .A1(n529), .A2(n514), .ZN(n407) );
  XNOR2_X1 U410 ( .A(n470), .B(n472), .ZN(n363) );
  XOR2_X1 U411 ( .A(G116), .B(KEYINPUT5), .Z(n489) );
  XOR2_X1 U412 ( .A(KEYINPUT12), .B(G122), .Z(n444) );
  XNOR2_X1 U413 ( .A(G113), .B(G104), .ZN(n443) );
  XOR2_X1 U414 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n447) );
  XNOR2_X1 U415 ( .A(G143), .B(G131), .ZN(n449) );
  XNOR2_X1 U416 ( .A(n458), .B(n438), .ZN(n704) );
  XNOR2_X1 U417 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n435) );
  XOR2_X1 U418 ( .A(G137), .B(G131), .Z(n436) );
  NAND2_X1 U419 ( .A1(n707), .A2(G227), .ZN(n396) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT97), .ZN(n394) );
  XNOR2_X1 U421 ( .A(n373), .B(n423), .ZN(n428) );
  XNOR2_X1 U422 ( .A(n697), .B(n422), .ZN(n373) );
  XNOR2_X1 U423 ( .A(n417), .B(KEYINPUT4), .ZN(n418) );
  XNOR2_X1 U424 ( .A(n569), .B(KEYINPUT107), .ZN(n359) );
  NAND2_X1 U425 ( .A1(n367), .A2(n350), .ZN(n529) );
  NOR2_X1 U426 ( .A1(n573), .A2(n368), .ZN(n367) );
  INV_X1 U427 ( .A(n513), .ZN(n368) );
  NOR2_X1 U428 ( .A1(n511), .A2(n507), .ZN(n521) );
  INV_X1 U429 ( .A(KEYINPUT22), .ZN(n364) );
  NAND2_X1 U430 ( .A1(n550), .A2(n485), .ZN(n388) );
  INV_X1 U431 ( .A(n527), .ZN(n522) );
  XNOR2_X1 U432 ( .A(n462), .B(n703), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U434 ( .A(n362), .B(n461), .ZN(n462) );
  XNOR2_X1 U435 ( .A(n386), .B(n384), .ZN(n686) );
  XNOR2_X1 U436 ( .A(n457), .B(n387), .ZN(n386) );
  XNOR2_X1 U437 ( .A(n458), .B(n385), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n454), .B(n453), .ZN(n387) );
  OR2_X1 U439 ( .A1(n539), .A2(n555), .ZN(n382) );
  INV_X1 U440 ( .A(KEYINPUT70), .ZN(n380) );
  INV_X1 U441 ( .A(KEYINPUT105), .ZN(n377) );
  XNOR2_X1 U442 ( .A(KEYINPUT15), .B(G902), .ZN(n579) );
  INV_X1 U443 ( .A(G469), .ZN(n398) );
  XNOR2_X1 U444 ( .A(n421), .B(G122), .ZN(n455) );
  XNOR2_X1 U445 ( .A(G116), .B(G107), .ZN(n421) );
  XOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n420) );
  NOR2_X1 U447 ( .A1(n630), .A2(n403), .ZN(n402) );
  INV_X1 U448 ( .A(n629), .ZN(n403) );
  NOR2_X1 U449 ( .A1(G902), .A2(G237), .ZN(n429) );
  AND2_X1 U450 ( .A1(n643), .A2(n486), .ZN(n504) );
  XNOR2_X1 U451 ( .A(n496), .B(n495), .ZN(n600) );
  XNOR2_X1 U452 ( .A(n492), .B(KEYINPUT16), .ZN(n409) );
  XNOR2_X1 U453 ( .A(n370), .B(n460), .ZN(n362) );
  XNOR2_X1 U454 ( .A(KEYINPUT83), .B(KEYINPUT72), .ZN(n460) );
  XNOR2_X1 U455 ( .A(n371), .B(KEYINPUT23), .ZN(n370) );
  INV_X1 U456 ( .A(KEYINPUT98), .ZN(n371) );
  XOR2_X1 U457 ( .A(KEYINPUT80), .B(KEYINPUT24), .Z(n461) );
  XNOR2_X1 U458 ( .A(G128), .B(G137), .ZN(n464) );
  XOR2_X1 U459 ( .A(G110), .B(G119), .Z(n465) );
  XOR2_X1 U460 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n454) );
  XNOR2_X1 U461 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n453) );
  INV_X1 U462 ( .A(n455), .ZN(n385) );
  XNOR2_X1 U463 ( .A(n452), .B(n451), .ZN(n592) );
  NAND2_X1 U464 ( .A1(G234), .A2(G237), .ZN(n473) );
  XOR2_X1 U465 ( .A(KEYINPUT94), .B(KEYINPUT14), .Z(n474) );
  INV_X1 U466 ( .A(KEYINPUT19), .ZN(n519) );
  NAND2_X1 U467 ( .A1(n512), .A2(n646), .ZN(n573) );
  XNOR2_X1 U468 ( .A(n496), .B(n440), .ZN(n681) );
  XOR2_X1 U469 ( .A(n427), .B(n426), .Z(n587) );
  XNOR2_X1 U470 ( .A(n510), .B(KEYINPUT42), .ZN(n720) );
  XNOR2_X1 U471 ( .A(n406), .B(KEYINPUT40), .ZN(n721) );
  XNOR2_X1 U472 ( .A(n562), .B(KEYINPUT35), .ZN(n716) );
  XNOR2_X1 U473 ( .A(n551), .B(KEYINPUT106), .ZN(n361) );
  XNOR2_X1 U474 ( .A(n688), .B(n689), .ZN(n366) );
  XNOR2_X1 U475 ( .A(n685), .B(n686), .ZN(n358) );
  INV_X1 U476 ( .A(n382), .ZN(n626) );
  XOR2_X1 U477 ( .A(n400), .B(n354), .Z(n350) );
  XOR2_X1 U478 ( .A(KEYINPUT13), .B(G475), .Z(n351) );
  AND2_X1 U479 ( .A1(n643), .A2(n649), .ZN(n352) );
  XNOR2_X1 U480 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n353) );
  XNOR2_X1 U481 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n354) );
  NAND2_X1 U482 ( .A1(n361), .A2(n352), .ZN(n613) );
  XOR2_X1 U483 ( .A(KEYINPUT64), .B(n516), .Z(n355) );
  XOR2_X1 U484 ( .A(n600), .B(n599), .Z(n356) );
  XOR2_X1 U485 ( .A(KEYINPUT65), .B(n580), .Z(n357) );
  NOR2_X2 U486 ( .A1(n606), .A2(n575), .ZN(n576) );
  NOR2_X2 U487 ( .A1(n643), .A2(n567), .ZN(n606) );
  NOR2_X1 U488 ( .A1(n358), .A2(n690), .ZN(G63) );
  NAND2_X1 U489 ( .A1(n359), .A2(n554), .ZN(n360) );
  XNOR2_X2 U490 ( .A(n360), .B(n353), .ZN(n667) );
  NOR2_X2 U491 ( .A1(n557), .A2(n388), .ZN(n365) );
  NAND2_X1 U492 ( .A1(n720), .A2(n721), .ZN(n517) );
  XNOR2_X2 U493 ( .A(n365), .B(n364), .ZN(n552) );
  NOR2_X1 U494 ( .A1(n366), .A2(n690), .ZN(G66) );
  XNOR2_X1 U495 ( .A(n468), .B(n369), .ZN(n689) );
  NAND2_X1 U496 ( .A1(n372), .A2(n357), .ZN(n585) );
  NAND2_X1 U497 ( .A1(n410), .A2(n414), .ZN(n372) );
  NOR2_X2 U498 ( .A1(n552), .A2(n554), .ZN(n564) );
  XNOR2_X1 U499 ( .A(n432), .B(n434), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n395), .B(n394), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n374), .B(KEYINPUT44), .ZN(n392) );
  NOR2_X1 U502 ( .A1(n552), .A2(n645), .ZN(n551) );
  NAND2_X1 U503 ( .A1(n541), .A2(n621), .ZN(n406) );
  NAND2_X1 U504 ( .A1(n405), .A2(n375), .ZN(n404) );
  XNOR2_X1 U505 ( .A(n517), .B(n355), .ZN(n375) );
  NAND2_X2 U506 ( .A1(n518), .A2(n658), .ZN(n535) );
  XNOR2_X1 U507 ( .A(n706), .B(KEYINPUT79), .ZN(n414) );
  XNOR2_X2 U508 ( .A(n583), .B(KEYINPUT86), .ZN(n706) );
  NAND2_X1 U509 ( .A1(n376), .A2(n402), .ZN(n583) );
  XNOR2_X1 U510 ( .A(n404), .B(n540), .ZN(n376) );
  INV_X1 U511 ( .A(n614), .ZN(n623) );
  INV_X1 U512 ( .A(n523), .ZN(n663) );
  XNOR2_X1 U513 ( .A(n378), .B(n377), .ZN(n523) );
  NAND2_X1 U514 ( .A1(n614), .A2(n379), .ZN(n378) );
  INV_X1 U515 ( .A(n621), .ZN(n379) );
  NAND2_X1 U516 ( .A1(n718), .A2(n613), .ZN(n393) );
  XNOR2_X2 U517 ( .A(n389), .B(KEYINPUT32), .ZN(n718) );
  NAND2_X1 U518 ( .A1(n564), .A2(n553), .ZN(n389) );
  NAND2_X1 U519 ( .A1(n576), .A2(n392), .ZN(n578) );
  INV_X4 U520 ( .A(G953), .ZN(n707) );
  XNOR2_X2 U521 ( .A(n399), .B(n397), .ZN(n511) );
  NAND2_X1 U522 ( .A1(n568), .A2(n658), .ZN(n400) );
  XNOR2_X2 U523 ( .A(n498), .B(n497), .ZN(n568) );
  XNOR2_X2 U524 ( .A(n401), .B(G143), .ZN(n437) );
  XNOR2_X2 U525 ( .A(n408), .B(G119), .ZN(n492) );
  XNOR2_X2 U526 ( .A(G113), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U527 ( .A(n412), .B(n411), .ZN(n410) );
  INV_X1 U528 ( .A(KEYINPUT85), .ZN(n411) );
  NOR2_X2 U529 ( .A1(n581), .A2(n579), .ZN(n412) );
  XNOR2_X2 U530 ( .A(n535), .B(n519), .ZN(n547) );
  XNOR2_X2 U531 ( .A(n431), .B(n413), .ZN(n518) );
  XNOR2_X1 U532 ( .A(n683), .B(n682), .ZN(n684) );
  AND2_X2 U533 ( .A1(n585), .A2(n584), .ZN(n679) );
  XNOR2_X2 U534 ( .A(n578), .B(n577), .ZN(n581) );
  INV_X1 U535 ( .A(KEYINPUT48), .ZN(n540) );
  XNOR2_X1 U536 ( .A(n416), .B(n696), .ZN(n432) );
  XNOR2_X1 U537 ( .A(n432), .B(n418), .ZN(n423) );
  INV_X1 U538 ( .A(KEYINPUT0), .ZN(n548) );
  INV_X1 U539 ( .A(KEYINPUT71), .ZN(n441) );
  XNOR2_X1 U540 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n604) );
  XNOR2_X1 U541 ( .A(n596), .B(KEYINPUT66), .ZN(n597) );
  XNOR2_X1 U542 ( .A(n491), .B(KEYINPUT73), .ZN(n416) );
  XNOR2_X1 U543 ( .A(n415), .B(KEYINPUT78), .ZN(n696) );
  XNOR2_X1 U544 ( .A(n437), .B(n442), .ZN(n417) );
  NAND2_X1 U545 ( .A1(G224), .A2(n707), .ZN(n419) );
  XOR2_X1 U546 ( .A(n420), .B(n419), .Z(n422) );
  BUF_X1 U547 ( .A(n428), .Z(n427) );
  XOR2_X1 U548 ( .A(KEYINPUT82), .B(KEYINPUT91), .Z(n425) );
  XNOR2_X1 U549 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n424) );
  XNOR2_X1 U550 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U551 ( .A1(n428), .A2(n579), .ZN(n431) );
  XNOR2_X1 U552 ( .A(n429), .B(KEYINPUT77), .ZN(n500) );
  NAND2_X1 U553 ( .A1(n500), .A2(G210), .ZN(n430) );
  XNOR2_X1 U554 ( .A(n433), .B(G107), .ZN(n434) );
  XNOR2_X1 U555 ( .A(n436), .B(n435), .ZN(n438) );
  INV_X1 U556 ( .A(n555), .ZN(n645) );
  XNOR2_X1 U557 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n703), .B(n445), .ZN(n452) );
  NAND2_X1 U559 ( .A1(G214), .A2(n487), .ZN(n446) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U561 ( .A(n448), .B(KEYINPUT101), .Z(n450) );
  XNOR2_X1 U562 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U563 ( .A1(G234), .A2(n707), .ZN(n456) );
  XOR2_X1 U564 ( .A(KEYINPUT8), .B(n456), .Z(n463) );
  NAND2_X1 U565 ( .A1(G217), .A2(n463), .ZN(n457) );
  NOR2_X1 U566 ( .A1(G902), .A2(n686), .ZN(n459) );
  XOR2_X1 U567 ( .A(G478), .B(n459), .Z(n526) );
  INV_X1 U568 ( .A(KEYINPUT25), .ZN(n472) );
  AND2_X1 U569 ( .A1(G221), .A2(n463), .ZN(n467) );
  XNOR2_X1 U570 ( .A(n465), .B(n464), .ZN(n466) );
  NOR2_X1 U571 ( .A1(G902), .A2(n689), .ZN(n471) );
  NAND2_X1 U572 ( .A1(n579), .A2(G234), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n469), .B(KEYINPUT20), .ZN(n482) );
  NAND2_X1 U574 ( .A1(G217), .A2(n482), .ZN(n470) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U576 ( .A(KEYINPUT76), .B(n475), .Z(n478) );
  AND2_X1 U577 ( .A1(G953), .A2(n478), .ZN(n476) );
  NAND2_X1 U578 ( .A1(G902), .A2(n476), .ZN(n542) );
  NOR2_X1 U579 ( .A1(G900), .A2(n542), .ZN(n477) );
  XNOR2_X1 U580 ( .A(n477), .B(KEYINPUT109), .ZN(n481) );
  NAND2_X1 U581 ( .A1(G952), .A2(n478), .ZN(n674) );
  NOR2_X1 U582 ( .A1(n674), .A2(G953), .ZN(n479) );
  XOR2_X1 U583 ( .A(n479), .B(KEYINPUT95), .Z(n545) );
  INV_X1 U584 ( .A(n545), .ZN(n480) );
  NAND2_X1 U585 ( .A1(n481), .A2(n480), .ZN(n513) );
  XOR2_X1 U586 ( .A(KEYINPUT21), .B(KEYINPUT99), .Z(n484) );
  NAND2_X1 U587 ( .A1(n482), .A2(G221), .ZN(n483) );
  XNOR2_X1 U588 ( .A(n484), .B(n483), .ZN(n642) );
  INV_X1 U589 ( .A(n642), .ZN(n485) );
  AND2_X1 U590 ( .A1(n513), .A2(n485), .ZN(n486) );
  NAND2_X1 U591 ( .A1(n487), .A2(G210), .ZN(n488) );
  XNOR2_X1 U592 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U593 ( .A(n490), .B(KEYINPUT100), .Z(n494) );
  XNOR2_X1 U594 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U596 ( .A1(n504), .A2(n554), .ZN(n499) );
  NOR2_X1 U597 ( .A1(n379), .A2(n499), .ZN(n534) );
  NAND2_X1 U598 ( .A1(G214), .A2(n500), .ZN(n658) );
  NAND2_X1 U599 ( .A1(n534), .A2(n658), .ZN(n501) );
  NOR2_X1 U600 ( .A1(n645), .A2(n501), .ZN(n502) );
  XNOR2_X1 U601 ( .A(n502), .B(KEYINPUT43), .ZN(n503) );
  NOR2_X1 U602 ( .A1(n532), .A2(n503), .ZN(n630) );
  INV_X1 U603 ( .A(KEYINPUT28), .ZN(n506) );
  AND2_X1 U604 ( .A1(n568), .A2(n504), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n507) );
  NAND2_X1 U606 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U607 ( .A1(n526), .A2(n527), .ZN(n550) );
  INV_X1 U608 ( .A(n550), .ZN(n661) );
  XNOR2_X1 U609 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n508) );
  XNOR2_X1 U610 ( .A(n509), .B(n508), .ZN(n655) );
  NAND2_X1 U611 ( .A1(n521), .A2(n655), .ZN(n510) );
  INV_X1 U612 ( .A(n659), .ZN(n514) );
  INV_X1 U613 ( .A(n511), .ZN(n512) );
  INV_X1 U614 ( .A(KEYINPUT39), .ZN(n515) );
  XOR2_X1 U615 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n516) );
  INV_X1 U616 ( .A(n547), .ZN(n520) );
  NAND2_X1 U617 ( .A1(n521), .A2(n520), .ZN(n619) );
  NAND2_X1 U618 ( .A1(n522), .A2(n526), .ZN(n614) );
  NAND2_X1 U619 ( .A1(KEYINPUT68), .A2(n523), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n525), .B(KEYINPUT47), .ZN(n533) );
  NAND2_X1 U621 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U622 ( .A(n528), .B(KEYINPUT108), .Z(n560) );
  INV_X1 U623 ( .A(n560), .ZN(n530) );
  NOR2_X1 U624 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U625 ( .A1(n532), .A2(n531), .ZN(n618) );
  XOR2_X1 U626 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n538) );
  INV_X1 U627 ( .A(n534), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U629 ( .A1(n623), .A2(n541), .ZN(n629) );
  NOR2_X1 U630 ( .A1(G898), .A2(n542), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n543), .B(KEYINPUT96), .ZN(n544) );
  NOR2_X1 U632 ( .A1(n545), .A2(n544), .ZN(n546) );
  AND2_X1 U633 ( .A1(n643), .A2(n645), .ZN(n553) );
  INV_X1 U634 ( .A(n555), .ZN(n556) );
  INV_X1 U635 ( .A(n557), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n667), .A2(n571), .ZN(n559) );
  XNOR2_X1 U637 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n558) );
  XNOR2_X1 U638 ( .A(n559), .B(n558), .ZN(n561) );
  NAND2_X1 U639 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U640 ( .A(KEYINPUT88), .ZN(n563) );
  XNOR2_X1 U641 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U642 ( .A(n566), .B(KEYINPUT89), .ZN(n567) );
  INV_X1 U643 ( .A(n568), .ZN(n649) );
  NOR2_X1 U644 ( .A1(n649), .A2(n569), .ZN(n653) );
  NAND2_X1 U645 ( .A1(n653), .A2(n571), .ZN(n570) );
  XNOR2_X1 U646 ( .A(KEYINPUT31), .B(n570), .ZN(n624) );
  NAND2_X1 U647 ( .A1(n649), .A2(n571), .ZN(n572) );
  NOR2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n609) );
  NOR2_X1 U649 ( .A1(n624), .A2(n609), .ZN(n574) );
  NOR2_X1 U650 ( .A1(n663), .A2(n574), .ZN(n575) );
  INV_X1 U651 ( .A(KEYINPUT45), .ZN(n577) );
  INV_X1 U652 ( .A(KEYINPUT2), .ZN(n634) );
  OR2_X1 U653 ( .A1(n579), .A2(n634), .ZN(n580) );
  INV_X1 U654 ( .A(n581), .ZN(n691) );
  NAND2_X1 U655 ( .A1(n691), .A2(KEYINPUT2), .ZN(n582) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n638) );
  INV_X1 U657 ( .A(n638), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n679), .A2(G210), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(n587), .ZN(n589) );
  NOR2_X1 U660 ( .A1(G952), .A2(n707), .ZN(n588) );
  XNOR2_X1 U661 ( .A(KEYINPUT92), .B(n588), .ZN(n690) );
  INV_X1 U662 ( .A(n690), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n589), .A2(n602), .ZN(n591) );
  INV_X1 U664 ( .A(KEYINPUT56), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n591), .B(n590), .ZN(G51) );
  NAND2_X1 U666 ( .A1(n349), .A2(G475), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT59), .ZN(n593) );
  XNOR2_X1 U668 ( .A(n594), .B(n593), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n595), .A2(n602), .ZN(n598) );
  INV_X1 U670 ( .A(KEYINPUT60), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n598), .B(n597), .ZN(G60) );
  NAND2_X1 U672 ( .A1(n679), .A2(G472), .ZN(n601) );
  XOR2_X1 U673 ( .A(KEYINPUT62), .B(KEYINPUT113), .Z(n599) );
  XNOR2_X1 U674 ( .A(n601), .B(n356), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(n604), .ZN(G57) );
  XOR2_X1 U677 ( .A(n606), .B(G101), .Z(n607) );
  XNOR2_X1 U678 ( .A(KEYINPUT114), .B(n607), .ZN(G3) );
  NAND2_X1 U679 ( .A1(n609), .A2(n621), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(G104), .ZN(G6) );
  XOR2_X1 U681 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n611) );
  NAND2_X1 U682 ( .A1(n609), .A2(n623), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U684 ( .A(G107), .B(n612), .ZN(G9) );
  XNOR2_X1 U685 ( .A(G110), .B(n613), .ZN(G12) );
  NOR2_X1 U686 ( .A1(n614), .A2(n619), .ZN(n616) );
  XNOR2_X1 U687 ( .A(G128), .B(KEYINPUT29), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(G30) );
  XOR2_X1 U689 ( .A(G143), .B(KEYINPUT115), .Z(n617) );
  XNOR2_X1 U690 ( .A(n618), .B(n617), .ZN(G45) );
  NOR2_X1 U691 ( .A1(n379), .A2(n619), .ZN(n620) );
  XOR2_X1 U692 ( .A(G146), .B(n620), .Z(G48) );
  NAND2_X1 U693 ( .A1(n624), .A2(n621), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n622), .B(G113), .ZN(G15) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n625), .B(G116), .ZN(G18) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT116), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT37), .ZN(n628) );
  XNOR2_X1 U699 ( .A(G125), .B(n628), .ZN(G27) );
  XNOR2_X1 U700 ( .A(G134), .B(n629), .ZN(G36) );
  XNOR2_X1 U701 ( .A(G140), .B(n630), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n631), .B(KEYINPUT117), .ZN(G42) );
  NAND2_X1 U703 ( .A1(n667), .A2(n655), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT122), .ZN(n641) );
  NAND2_X1 U705 ( .A1(n634), .A2(n706), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n633), .B(KEYINPUT84), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n634), .A2(n581), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U710 ( .A1(G953), .A2(n639), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n677) );
  XNOR2_X1 U712 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n673) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n644), .B(KEYINPUT49), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT50), .B(n647), .Z(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U720 ( .A(KEYINPUT51), .B(n654), .ZN(n656) );
  NAND2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n657), .B(KEYINPUT118), .ZN(n670) );
  NOR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U726 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U727 ( .A(n666), .B(KEYINPUT119), .ZN(n668) );
  NAND2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U730 ( .A(n671), .B(KEYINPUT52), .ZN(n672) );
  XNOR2_X1 U731 ( .A(n673), .B(n672), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U734 ( .A(KEYINPUT53), .B(n678), .ZN(G75) );
  BUF_X2 U735 ( .A(n349), .Z(n687) );
  NAND2_X1 U736 ( .A1(n687), .A2(G469), .ZN(n683) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n680) );
  XNOR2_X1 U738 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U739 ( .A1(n690), .A2(n684), .ZN(G54) );
  NAND2_X1 U740 ( .A1(G478), .A2(n687), .ZN(n685) );
  NAND2_X1 U741 ( .A1(G217), .A2(n687), .ZN(n688) );
  NAND2_X1 U742 ( .A1(n707), .A2(n691), .ZN(n695) );
  NAND2_X1 U743 ( .A1(G953), .A2(G224), .ZN(n692) );
  XNOR2_X1 U744 ( .A(KEYINPUT61), .B(n692), .ZN(n693) );
  NAND2_X1 U745 ( .A1(n693), .A2(G898), .ZN(n694) );
  NAND2_X1 U746 ( .A1(n695), .A2(n694), .ZN(n702) );
  XNOR2_X1 U747 ( .A(G101), .B(n696), .ZN(n698) );
  XNOR2_X1 U748 ( .A(n698), .B(n697), .ZN(n700) );
  NOR2_X1 U749 ( .A1(G898), .A2(n707), .ZN(n699) );
  NOR2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U751 ( .A(n702), .B(n701), .ZN(G69) );
  XNOR2_X1 U752 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U753 ( .A(n705), .B(KEYINPUT123), .ZN(n709) );
  XOR2_X1 U754 ( .A(n706), .B(n709), .Z(n708) );
  NAND2_X1 U755 ( .A1(n708), .A2(n707), .ZN(n714) );
  XNOR2_X1 U756 ( .A(G227), .B(n709), .ZN(n710) );
  NAND2_X1 U757 ( .A1(n710), .A2(G900), .ZN(n711) );
  XOR2_X1 U758 ( .A(KEYINPUT124), .B(n711), .Z(n712) );
  NAND2_X1 U759 ( .A1(n712), .A2(G953), .ZN(n713) );
  NAND2_X1 U760 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U761 ( .A(KEYINPUT125), .B(n715), .ZN(G72) );
  XOR2_X1 U762 ( .A(n716), .B(G122), .Z(n717) );
  XNOR2_X1 U763 ( .A(KEYINPUT126), .B(n717), .ZN(G24) );
  XOR2_X1 U764 ( .A(n718), .B(G119), .Z(n719) );
  XNOR2_X1 U765 ( .A(KEYINPUT127), .B(n719), .ZN(G21) );
  XNOR2_X1 U766 ( .A(n720), .B(G137), .ZN(G39) );
  XNOR2_X1 U767 ( .A(G131), .B(n721), .ZN(G33) );
endmodule

