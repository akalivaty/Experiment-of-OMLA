

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719;

  XNOR2_X1 U366 ( .A(n425), .B(KEYINPUT65), .ZN(n424) );
  NAND2_X1 U367 ( .A1(n630), .A2(n707), .ZN(n383) );
  XNOR2_X2 U368 ( .A(G125), .B(G146), .ZN(n437) );
  XNOR2_X2 U369 ( .A(n388), .B(KEYINPUT22), .ZN(n519) );
  XNOR2_X2 U370 ( .A(n597), .B(n596), .ZN(n599) );
  OR2_X2 U371 ( .A1(n536), .A2(n389), .ZN(n388) );
  NOR2_X1 U372 ( .A1(n521), .A2(n645), .ZN(n535) );
  XNOR2_X1 U373 ( .A(n418), .B(n417), .ZN(n536) );
  NOR2_X1 U374 ( .A1(n561), .A2(n484), .ZN(n418) );
  XNOR2_X1 U375 ( .A(n477), .B(n476), .ZN(n590) );
  NOR2_X1 U376 ( .A1(n640), .A2(n639), .ZN(n376) );
  XNOR2_X1 U377 ( .A(n573), .B(n572), .ZN(n640) );
  OR2_X1 U378 ( .A1(n639), .A2(n390), .ZN(n389) );
  INV_X1 U379 ( .A(n590), .ZN(n580) );
  XNOR2_X1 U380 ( .A(n460), .B(G134), .ZN(n498) );
  XNOR2_X1 U381 ( .A(n361), .B(G101), .ZN(n500) );
  XNOR2_X1 U382 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U383 ( .A(n423), .B(n422), .ZN(n717) );
  NOR2_X1 U384 ( .A1(G902), .A2(G237), .ZN(n456) );
  NOR2_X1 U385 ( .A1(n717), .A2(n349), .ZN(n396) );
  XOR2_X1 U386 ( .A(G140), .B(KEYINPUT69), .Z(n499) );
  NOR2_X1 U387 ( .A1(G902), .A2(n679), .ZN(n444) );
  XNOR2_X1 U388 ( .A(n449), .B(n450), .ZN(n490) );
  XOR2_X1 U389 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n450) );
  XNOR2_X1 U390 ( .A(KEYINPUT10), .B(n437), .ZN(n700) );
  XNOR2_X1 U391 ( .A(n523), .B(n522), .ZN(n667) );
  XNOR2_X1 U392 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n522) );
  XNOR2_X1 U393 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U394 ( .A1(n683), .A2(G217), .ZN(n401) );
  XNOR2_X1 U395 ( .A(n511), .B(n509), .ZN(n413) );
  NOR2_X1 U396 ( .A1(n641), .A2(n620), .ZN(n562) );
  INV_X1 U397 ( .A(n619), .ZN(n570) );
  NAND2_X1 U398 ( .A1(n395), .A2(n396), .ZN(n394) );
  AND2_X1 U399 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U400 ( .A(n498), .B(n497), .ZN(n508) );
  XNOR2_X1 U401 ( .A(KEYINPUT4), .B(G131), .ZN(n496) );
  INV_X1 U402 ( .A(KEYINPUT67), .ZN(n361) );
  NAND2_X1 U403 ( .A1(n653), .A2(n636), .ZN(n416) );
  XNOR2_X1 U404 ( .A(KEYINPUT70), .B(n556), .ZN(n578) );
  XNOR2_X1 U405 ( .A(n506), .B(n505), .ZN(n559) );
  INV_X1 U406 ( .A(G469), .ZN(n505) );
  XNOR2_X1 U407 ( .A(n419), .B(n469), .ZN(n512) );
  XNOR2_X1 U408 ( .A(n421), .B(n420), .ZN(n419) );
  INV_X1 U409 ( .A(G119), .ZN(n420) );
  XNOR2_X1 U410 ( .A(G104), .B(G110), .ZN(n467) );
  XNOR2_X1 U411 ( .A(KEYINPUT16), .B(G122), .ZN(n364) );
  XOR2_X1 U412 ( .A(G143), .B(G122), .Z(n436) );
  XNOR2_X1 U413 ( .A(G113), .B(G104), .ZN(n435) );
  XNOR2_X1 U414 ( .A(n443), .B(KEYINPUT96), .ZN(n408) );
  XNOR2_X1 U415 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U416 ( .A(G140), .B(G131), .ZN(n438) );
  XNOR2_X1 U417 ( .A(n376), .B(n347), .ZN(n666) );
  XNOR2_X1 U418 ( .A(n411), .B(n410), .ZN(n592) );
  INV_X1 U419 ( .A(KEYINPUT39), .ZN(n410) );
  NOR2_X1 U420 ( .A1(n536), .A2(n667), .ZN(n525) );
  INV_X1 U421 ( .A(n649), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n384), .B(n344), .ZN(n561) );
  NAND2_X1 U423 ( .A1(n542), .A2(n557), .ZN(n425) );
  INV_X1 U424 ( .A(n538), .ZN(n539) );
  XNOR2_X1 U425 ( .A(n517), .B(KEYINPUT101), .ZN(n577) );
  XNOR2_X1 U426 ( .A(n493), .B(n700), .ZN(n684) );
  XNOR2_X1 U427 ( .A(n383), .B(n631), .ZN(n598) );
  NAND2_X1 U428 ( .A1(n424), .A2(n555), .ZN(n395) );
  NAND2_X1 U429 ( .A1(G234), .A2(G237), .ZN(n479) );
  XNOR2_X1 U430 ( .A(n412), .B(n359), .ZN(n600) );
  XNOR2_X1 U431 ( .A(n360), .B(n514), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n413), .B(n508), .ZN(n412) );
  XNOR2_X1 U433 ( .A(n403), .B(KEYINPUT73), .ZN(n402) );
  INV_X1 U434 ( .A(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U435 ( .A(G116), .B(G107), .ZN(n446) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT75), .ZN(n510) );
  NAND2_X1 U437 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U438 ( .A(G237), .ZN(n371) );
  XOR2_X1 U439 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n439) );
  XNOR2_X1 U440 ( .A(n500), .B(n457), .ZN(n459) );
  INV_X1 U441 ( .A(n520), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n495), .B(KEYINPUT25), .ZN(n381) );
  XNOR2_X1 U443 ( .A(G119), .B(G137), .ZN(n485) );
  XOR2_X1 U444 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n487) );
  AND2_X1 U445 ( .A1(n373), .A2(n577), .ZN(n579) );
  NOR2_X1 U446 ( .A1(n578), .A2(n624), .ZN(n373) );
  NOR2_X1 U447 ( .A1(n580), .A2(n586), .ZN(n582) );
  NOR2_X1 U448 ( .A1(n567), .A2(n566), .ZN(n571) );
  INV_X1 U449 ( .A(n565), .ZN(n414) );
  XNOR2_X1 U450 ( .A(n416), .B(n564), .ZN(n415) );
  INV_X1 U451 ( .A(KEYINPUT0), .ZN(n417) );
  INV_X1 U452 ( .A(n653), .ZN(n557) );
  INV_X1 U453 ( .A(KEYINPUT64), .ZN(n380) );
  XNOR2_X1 U454 ( .A(n364), .B(n363), .ZN(n468) );
  INV_X1 U455 ( .A(KEYINPUT72), .ZN(n363) );
  XNOR2_X1 U456 ( .A(n407), .B(n406), .ZN(n679) );
  XNOR2_X1 U457 ( .A(n343), .B(n700), .ZN(n406) );
  XNOR2_X1 U458 ( .A(n442), .B(n408), .ZN(n407) );
  INV_X1 U459 ( .A(G953), .ZN(n372) );
  NAND2_X1 U460 ( .A1(n345), .A2(n668), .ZN(n354) );
  XNOR2_X1 U461 ( .A(n409), .B(n348), .ZN(n715) );
  NOR2_X1 U462 ( .A1(n592), .A2(n624), .ZN(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT32), .B(KEYINPUT80), .ZN(n422) );
  NOR2_X1 U464 ( .A1(n519), .A2(n365), .ZN(n423) );
  NAND2_X1 U465 ( .A1(n518), .A2(n366), .ZN(n365) );
  NAND2_X1 U466 ( .A1(n368), .A2(n367), .ZN(n620) );
  INV_X1 U467 ( .A(n561), .ZN(n367) );
  INV_X1 U468 ( .A(n574), .ZN(n368) );
  NAND2_X1 U469 ( .A1(n399), .A2(n357), .ZN(n398) );
  XNOR2_X1 U470 ( .A(n401), .B(n400), .ZN(n399) );
  INV_X1 U471 ( .A(KEYINPUT120), .ZN(n355) );
  XNOR2_X1 U472 ( .A(n427), .B(n426), .ZN(G75) );
  INV_X1 U473 ( .A(KEYINPUT53), .ZN(n426) );
  NAND2_X1 U474 ( .A1(n428), .A2(n372), .ZN(n427) );
  XNOR2_X1 U475 ( .A(n429), .B(KEYINPUT117), .ZN(n428) );
  INV_X1 U476 ( .A(n395), .ZN(n615) );
  XNOR2_X1 U477 ( .A(n382), .B(n381), .ZN(n549) );
  AND2_X1 U478 ( .A1(n555), .A2(n349), .ZN(n342) );
  XOR2_X1 U479 ( .A(n436), .B(n435), .Z(n343) );
  XOR2_X1 U480 ( .A(n478), .B(KEYINPUT76), .Z(n344) );
  OR2_X1 U481 ( .A1(n664), .A2(n663), .ZN(n345) );
  OR2_X1 U482 ( .A1(n383), .A2(n631), .ZN(n346) );
  NAND2_X1 U483 ( .A1(n540), .A2(n539), .ZN(n624) );
  XNOR2_X1 U484 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n347) );
  XNOR2_X1 U485 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n348) );
  AND2_X1 U486 ( .A1(n530), .A2(KEYINPUT84), .ZN(n349) );
  NOR2_X1 U487 ( .A1(n708), .A2(G952), .ZN(n685) );
  INV_X1 U488 ( .A(n685), .ZN(n357) );
  XOR2_X1 U489 ( .A(n602), .B(n601), .Z(n350) );
  XNOR2_X1 U490 ( .A(n679), .B(KEYINPUT59), .ZN(n351) );
  XNOR2_X1 U491 ( .A(n672), .B(n671), .ZN(n352) );
  XOR2_X1 U492 ( .A(KEYINPUT118), .B(KEYINPUT56), .Z(n353) );
  NAND2_X1 U493 ( .A1(n590), .A2(n636), .ZN(n384) );
  NAND2_X1 U494 ( .A1(n394), .A2(n391), .ZN(n397) );
  XNOR2_X1 U495 ( .A(n385), .B(n353), .ZN(G51) );
  XNOR2_X1 U496 ( .A(n460), .B(KEYINPUT4), .ZN(n464) );
  OR2_X1 U497 ( .A1(n665), .A2(n354), .ZN(n429) );
  XNOR2_X1 U498 ( .A(n356), .B(n355), .ZN(G63) );
  NAND2_X1 U499 ( .A1(n377), .A2(n357), .ZN(n356) );
  XNOR2_X1 U500 ( .A(n387), .B(n352), .ZN(n386) );
  NAND2_X1 U501 ( .A1(n386), .A2(n357), .ZN(n385) );
  AND2_X2 U502 ( .A1(n358), .A2(n357), .ZN(n369) );
  XNOR2_X1 U503 ( .A(n603), .B(n350), .ZN(n358) );
  NAND2_X1 U504 ( .A1(n415), .A2(n414), .ZN(n566) );
  INV_X1 U505 ( .A(n513), .ZN(n360) );
  AND2_X2 U506 ( .A1(n362), .A2(n357), .ZN(n681) );
  XNOR2_X1 U507 ( .A(n680), .B(n351), .ZN(n362) );
  NOR2_X1 U508 ( .A1(n600), .A2(G902), .ZN(n516) );
  XNOR2_X2 U509 ( .A(G143), .B(G128), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n375), .B(n374), .ZN(n595) );
  NAND2_X1 U511 ( .A1(n560), .A2(n559), .ZN(n574) );
  NOR2_X1 U512 ( .A1(n684), .A2(G902), .ZN(n382) );
  NAND2_X1 U513 ( .A1(n405), .A2(n402), .ZN(n375) );
  XNOR2_X1 U514 ( .A(n369), .B(n605), .ZN(G57) );
  XNOR2_X1 U515 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U516 ( .A(n682), .ZN(n378) );
  NAND2_X1 U517 ( .A1(n683), .A2(G478), .ZN(n379) );
  NOR2_X4 U518 ( .A1(n599), .A2(n598), .ZN(n683) );
  XNOR2_X2 U519 ( .A(n380), .B(G953), .ZN(n708) );
  NAND2_X1 U520 ( .A1(n383), .A2(KEYINPUT83), .ZN(n597) );
  NAND2_X1 U521 ( .A1(n683), .A2(G210), .ZN(n387) );
  NOR2_X2 U522 ( .A1(n519), .A2(n587), .ZN(n542) );
  NAND2_X1 U523 ( .A1(n717), .A2(n349), .ZN(n393) );
  NAND2_X1 U524 ( .A1(n424), .A2(n342), .ZN(n392) );
  NAND2_X1 U525 ( .A1(n397), .A2(n714), .ZN(n532) );
  XNOR2_X1 U526 ( .A(n398), .B(KEYINPUT121), .ZN(G66) );
  INV_X1 U527 ( .A(n684), .ZN(n400) );
  NAND2_X1 U528 ( .A1(n404), .A2(n570), .ZN(n403) );
  XNOR2_X1 U529 ( .A(n562), .B(KEYINPUT47), .ZN(n404) );
  AND2_X1 U530 ( .A1(n585), .A2(n713), .ZN(n405) );
  INV_X1 U531 ( .A(n437), .ZN(n457) );
  NOR2_X1 U532 ( .A1(n715), .A2(n719), .ZN(n576) );
  XNOR2_X2 U533 ( .A(n580), .B(KEYINPUT38), .ZN(n637) );
  XNOR2_X1 U534 ( .A(n463), .B(n464), .ZN(n465) );
  XNOR2_X1 U535 ( .A(n459), .B(n458), .ZN(n466) );
  NAND2_X1 U536 ( .A1(n571), .A2(n637), .ZN(n411) );
  XNOR2_X2 U537 ( .A(n516), .B(n515), .ZN(n653) );
  XNOR2_X1 U538 ( .A(n466), .B(n465), .ZN(n471) );
  AND2_X1 U539 ( .A1(G227), .A2(n708), .ZN(n430) );
  INV_X1 U540 ( .A(KEYINPUT97), .ZN(n440) );
  XNOR2_X1 U541 ( .A(n496), .B(G137), .ZN(n497) );
  INV_X1 U542 ( .A(KEYINPUT107), .ZN(n572) );
  XNOR2_X1 U543 ( .A(n468), .B(n502), .ZN(n470) );
  XNOR2_X1 U544 ( .A(n701), .B(n501), .ZN(n504) );
  INV_X1 U545 ( .A(KEYINPUT91), .ZN(n474) );
  INV_X1 U546 ( .A(G472), .ZN(n515) );
  AND2_X1 U547 ( .A1(n718), .A2(n593), .ZN(n594) );
  XNOR2_X1 U548 ( .A(n559), .B(n507), .ZN(n521) );
  XNOR2_X1 U549 ( .A(n604), .B(KEYINPUT88), .ZN(n605) );
  XOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .Z(n472) );
  INV_X1 U551 ( .A(n472), .ZN(n596) );
  NAND2_X1 U552 ( .A1(n596), .A2(G234), .ZN(n431) );
  XNOR2_X1 U553 ( .A(n431), .B(KEYINPUT20), .ZN(n494) );
  NAND2_X1 U554 ( .A1(G221), .A2(n494), .ZN(n432) );
  XNOR2_X1 U555 ( .A(KEYINPUT21), .B(n432), .ZN(n648) );
  XNOR2_X1 U556 ( .A(n648), .B(KEYINPUT95), .ZN(n520) );
  XOR2_X1 U557 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n434) );
  XNOR2_X1 U558 ( .A(KEYINPUT98), .B(G475), .ZN(n433) );
  XNOR2_X1 U559 ( .A(n434), .B(n433), .ZN(n445) );
  XNOR2_X1 U560 ( .A(n439), .B(n438), .ZN(n441) );
  NAND2_X1 U561 ( .A1(n510), .A2(G214), .ZN(n443) );
  XOR2_X1 U562 ( .A(n445), .B(n444), .Z(n538) );
  XOR2_X1 U563 ( .A(KEYINPUT9), .B(G122), .Z(n447) );
  XNOR2_X1 U564 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U565 ( .A(n498), .B(n448), .ZN(n454) );
  XOR2_X1 U566 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n452) );
  NAND2_X1 U567 ( .A1(G234), .A2(n708), .ZN(n449) );
  NAND2_X1 U568 ( .A1(G217), .A2(n490), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U570 ( .A(n454), .B(n453), .ZN(n682) );
  NOR2_X1 U571 ( .A1(G902), .A2(n682), .ZN(n455) );
  XNOR2_X1 U572 ( .A(G478), .B(n455), .ZN(n540) );
  NAND2_X1 U573 ( .A1(n538), .A2(n540), .ZN(n639) );
  XOR2_X1 U574 ( .A(KEYINPUT74), .B(n456), .Z(n473) );
  NAND2_X1 U575 ( .A1(n473), .A2(G214), .ZN(n636) );
  NAND2_X1 U576 ( .A1(G224), .A2(n708), .ZN(n458) );
  XOR2_X1 U577 ( .A(KEYINPUT18), .B(KEYINPUT90), .Z(n462) );
  XNOR2_X1 U578 ( .A(KEYINPUT77), .B(KEYINPUT17), .ZN(n461) );
  XNOR2_X1 U579 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U580 ( .A(n467), .B(G107), .ZN(n502) );
  XNOR2_X1 U581 ( .A(G116), .B(G113), .ZN(n469) );
  XNOR2_X1 U582 ( .A(n512), .B(n470), .ZN(n686) );
  XNOR2_X1 U583 ( .A(n471), .B(n686), .ZN(n672) );
  NOR2_X1 U584 ( .A1(n672), .A2(n472), .ZN(n477) );
  NAND2_X1 U585 ( .A1(n473), .A2(G210), .ZN(n475) );
  XNOR2_X1 U586 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n478) );
  XNOR2_X1 U587 ( .A(n479), .B(KEYINPUT14), .ZN(n480) );
  NAND2_X1 U588 ( .A1(n480), .A2(G952), .ZN(n664) );
  NOR2_X1 U589 ( .A1(G953), .A2(n664), .ZN(n553) );
  NAND2_X1 U590 ( .A1(G902), .A2(n480), .ZN(n550) );
  XOR2_X1 U591 ( .A(G898), .B(KEYINPUT92), .Z(n693) );
  NAND2_X1 U592 ( .A1(n693), .A2(G953), .ZN(n481) );
  XOR2_X1 U593 ( .A(KEYINPUT93), .B(n481), .Z(n687) );
  NOR2_X1 U594 ( .A1(n550), .A2(n687), .ZN(n482) );
  NOR2_X1 U595 ( .A1(n553), .A2(n482), .ZN(n483) );
  XNOR2_X1 U596 ( .A(n483), .B(KEYINPUT94), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n499), .B(n485), .ZN(n489) );
  XNOR2_X1 U598 ( .A(G110), .B(G128), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U600 ( .A(n489), .B(n488), .Z(n492) );
  NAND2_X1 U601 ( .A1(G221), .A2(n490), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U603 ( .A1(n494), .A2(G217), .ZN(n495) );
  XNOR2_X1 U604 ( .A(KEYINPUT102), .B(n549), .ZN(n649) );
  XNOR2_X1 U605 ( .A(n499), .B(n508), .ZN(n701) );
  XOR2_X1 U606 ( .A(n500), .B(G146), .Z(n513) );
  XNOR2_X1 U607 ( .A(n513), .B(n430), .ZN(n501) );
  INV_X1 U608 ( .A(n502), .ZN(n503) );
  XNOR2_X1 U609 ( .A(n504), .B(n503), .ZN(n673) );
  NOR2_X1 U610 ( .A1(n673), .A2(G902), .ZN(n506) );
  INV_X1 U611 ( .A(KEYINPUT1), .ZN(n507) );
  BUF_X1 U612 ( .A(n521), .Z(n646) );
  INV_X1 U613 ( .A(KEYINPUT5), .ZN(n509) );
  NAND2_X1 U614 ( .A1(n510), .A2(G210), .ZN(n511) );
  INV_X1 U615 ( .A(n512), .ZN(n514) );
  XNOR2_X1 U616 ( .A(n653), .B(KEYINPUT6), .ZN(n517) );
  NOR2_X1 U617 ( .A1(n646), .A2(n577), .ZN(n518) );
  INV_X1 U618 ( .A(n646), .ZN(n587) );
  INV_X1 U619 ( .A(KEYINPUT44), .ZN(n530) );
  NAND2_X1 U620 ( .A1(n549), .A2(n520), .ZN(n645) );
  NAND2_X1 U621 ( .A1(n535), .A2(n577), .ZN(n523) );
  XNOR2_X1 U622 ( .A(KEYINPUT34), .B(KEYINPUT79), .ZN(n524) );
  XNOR2_X1 U623 ( .A(n525), .B(n524), .ZN(n527) );
  NOR2_X1 U624 ( .A1(n538), .A2(n540), .ZN(n568) );
  XOR2_X1 U625 ( .A(n568), .B(KEYINPUT78), .Z(n526) );
  NOR2_X1 U626 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U627 ( .A(n528), .B(KEYINPUT35), .ZN(n714) );
  INV_X1 U628 ( .A(n714), .ZN(n529) );
  NAND2_X1 U629 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U630 ( .A1(n532), .A2(n531), .ZN(n546) );
  INV_X1 U631 ( .A(n645), .ZN(n533) );
  NAND2_X1 U632 ( .A1(n559), .A2(n533), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n536), .A2(n567), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n534), .A2(n557), .ZN(n609) );
  NAND2_X1 U635 ( .A1(n653), .A2(n535), .ZN(n656) );
  NOR2_X1 U636 ( .A1(n656), .A2(n536), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n537), .B(KEYINPUT31), .ZN(n626) );
  NAND2_X1 U638 ( .A1(n609), .A2(n626), .ZN(n541) );
  OR2_X1 U639 ( .A1(n540), .A2(n539), .ZN(n627) );
  NAND2_X1 U640 ( .A1(n624), .A2(n627), .ZN(n548) );
  AND2_X1 U641 ( .A1(n541), .A2(n548), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n649), .A2(n542), .ZN(n543) );
  NOR2_X1 U643 ( .A1(n577), .A2(n543), .ZN(n606) );
  NOR2_X1 U644 ( .A1(n544), .A2(n606), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X2 U646 ( .A(n547), .B(KEYINPUT45), .ZN(n630) );
  INV_X1 U647 ( .A(n548), .ZN(n641) );
  INV_X1 U648 ( .A(n549), .ZN(n555) );
  OR2_X1 U649 ( .A1(n708), .A2(n550), .ZN(n551) );
  NOR2_X1 U650 ( .A1(G900), .A2(n551), .ZN(n552) );
  NOR2_X1 U651 ( .A1(n553), .A2(n552), .ZN(n565) );
  NOR2_X1 U652 ( .A1(n565), .A2(n648), .ZN(n554) );
  NAND2_X1 U653 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U654 ( .A1(n578), .A2(n557), .ZN(n558) );
  XNOR2_X1 U655 ( .A(n558), .B(KEYINPUT28), .ZN(n560) );
  XNOR2_X1 U656 ( .A(KEYINPUT105), .B(KEYINPUT30), .ZN(n563) );
  XNOR2_X1 U657 ( .A(n563), .B(KEYINPUT104), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n571), .A2(n568), .ZN(n569) );
  NOR2_X1 U659 ( .A1(n580), .A2(n569), .ZN(n619) );
  NAND2_X1 U660 ( .A1(n637), .A2(n636), .ZN(n573) );
  NOR2_X1 U661 ( .A1(n574), .A2(n666), .ZN(n575) );
  XNOR2_X1 U662 ( .A(n575), .B(KEYINPUT42), .ZN(n719) );
  XNOR2_X1 U663 ( .A(n576), .B(KEYINPUT46), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n579), .A2(n636), .ZN(n586) );
  XNOR2_X1 U665 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n581) );
  XNOR2_X1 U666 ( .A(n582), .B(n581), .ZN(n583) );
  NOR2_X1 U667 ( .A1(n583), .A2(n646), .ZN(n584) );
  XNOR2_X1 U668 ( .A(n584), .B(KEYINPUT109), .ZN(n713) );
  NOR2_X1 U669 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U670 ( .A(n588), .B(KEYINPUT43), .ZN(n589) );
  NOR2_X1 U671 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U672 ( .A(KEYINPUT103), .B(n591), .ZN(n718) );
  NOR2_X1 U673 ( .A1(n592), .A2(n627), .ZN(n629) );
  INV_X1 U674 ( .A(n629), .ZN(n593) );
  AND2_X2 U675 ( .A1(n595), .A2(n594), .ZN(n707) );
  INV_X1 U676 ( .A(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U677 ( .A1(n683), .A2(G472), .ZN(n603) );
  XOR2_X1 U678 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n602) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT110), .ZN(n601) );
  INV_X1 U680 ( .A(KEYINPUT63), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n606), .B(G101), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT111), .ZN(G3) );
  NOR2_X1 U683 ( .A1(n624), .A2(n609), .ZN(n608) );
  XOR2_X1 U684 ( .A(G104), .B(n608), .Z(G6) );
  NOR2_X1 U685 ( .A1(n627), .A2(n609), .ZN(n614) );
  XOR2_X1 U686 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n611) );
  XNOR2_X1 U687 ( .A(G107), .B(KEYINPUT26), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U689 ( .A(KEYINPUT112), .B(n612), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n614), .B(n613), .ZN(G9) );
  XOR2_X1 U691 ( .A(G110), .B(n615), .Z(G12) );
  NOR2_X1 U692 ( .A1(n627), .A2(n620), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(G128), .B(n618), .ZN(G30) );
  XOR2_X1 U696 ( .A(G143), .B(n619), .Z(G45) );
  NOR2_X1 U697 ( .A1(n624), .A2(n620), .ZN(n622) );
  XNOR2_X1 U698 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U700 ( .A(G146), .B(n623), .ZN(G48) );
  NOR2_X1 U701 ( .A1(n624), .A2(n626), .ZN(n625) );
  XOR2_X1 U702 ( .A(G113), .B(n625), .Z(G15) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U704 ( .A(G116), .B(n628), .Z(G18) );
  XOR2_X1 U705 ( .A(G134), .B(n629), .Z(G36) );
  INV_X1 U706 ( .A(n630), .ZN(n694) );
  NAND2_X1 U707 ( .A1(n694), .A2(n631), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT82), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n346), .A2(n633), .ZN(n635) );
  NOR2_X1 U710 ( .A1(n707), .A2(KEYINPUT2), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n665) );
  NOR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n667), .A2(n644), .ZN(n661) );
  NAND2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(KEYINPUT50), .B(n647), .ZN(n655) );
  INV_X1 U719 ( .A(n648), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT49), .B(n651), .Z(n652) );
  NOR2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U725 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n666), .A2(n659), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(KEYINPUT52), .ZN(n663) );
  OR2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT81), .B(KEYINPUT86), .Z(n670) );
  XNOR2_X1 U731 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n669) );
  XNOR2_X1 U732 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U733 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n675) );
  XNOR2_X1 U734 ( .A(n673), .B(KEYINPUT119), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n675), .B(n674), .ZN(n677) );
  NAND2_X1 U736 ( .A1(n683), .A2(G469), .ZN(n676) );
  XOR2_X1 U737 ( .A(n677), .B(n676), .Z(n678) );
  NOR2_X1 U738 ( .A1(n685), .A2(n678), .ZN(G54) );
  NAND2_X1 U739 ( .A1(n683), .A2(G475), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n681), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U741 ( .A(n686), .B(G101), .ZN(n688) );
  NAND2_X1 U742 ( .A1(n688), .A2(n687), .ZN(n699) );
  XOR2_X1 U743 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n690) );
  NAND2_X1 U744 ( .A1(G224), .A2(G953), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n690), .B(n689), .ZN(n691) );
  XOR2_X1 U746 ( .A(KEYINPUT122), .B(n691), .Z(n692) );
  NOR2_X1 U747 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U748 ( .A1(G953), .A2(n694), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n695), .B(KEYINPUT124), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U751 ( .A(n699), .B(n698), .ZN(G69) );
  XOR2_X1 U752 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n703) );
  XNOR2_X1 U753 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U754 ( .A(n703), .B(n702), .ZN(n706) );
  XOR2_X1 U755 ( .A(G227), .B(n706), .Z(n704) );
  NAND2_X1 U756 ( .A1(G900), .A2(n704), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(G953), .ZN(n711) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U759 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U760 ( .A1(n711), .A2(n710), .ZN(G72) );
  XOR2_X1 U761 ( .A(G125), .B(KEYINPUT37), .Z(n712) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(G27) );
  XNOR2_X1 U763 ( .A(G122), .B(n714), .ZN(G24) );
  XNOR2_X1 U764 ( .A(n715), .B(G131), .ZN(n716) );
  XNOR2_X1 U765 ( .A(n716), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U766 ( .A(n717), .B(G119), .Z(G21) );
  XNOR2_X1 U767 ( .A(G140), .B(n718), .ZN(G42) );
  XOR2_X1 U768 ( .A(G137), .B(n719), .Z(G39) );
endmodule

