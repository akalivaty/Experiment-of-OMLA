

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U323 ( .A(n547), .B(KEYINPUT123), .ZN(n548) );
  NOR2_X1 U324 ( .A1(n555), .A2(n554), .ZN(n566) );
  XOR2_X1 U325 ( .A(G190GAT), .B(G99GAT), .Z(n291) );
  XOR2_X1 U326 ( .A(n408), .B(n316), .Z(n292) );
  XNOR2_X1 U327 ( .A(n417), .B(n416), .ZN(n581) );
  XNOR2_X1 U328 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U329 ( .A(n404), .B(n403), .ZN(n406) );
  NOR2_X1 U330 ( .A1(n550), .A2(n518), .ZN(n327) );
  OR2_X1 U331 ( .A1(n585), .A2(n581), .ZN(n418) );
  XNOR2_X1 U332 ( .A(n549), .B(n548), .ZN(n570) );
  XOR2_X1 U333 ( .A(KEYINPUT96), .B(n328), .Z(n571) );
  XNOR2_X1 U334 ( .A(n415), .B(n414), .ZN(n416) );
  AND2_X1 U335 ( .A1(n492), .A2(n457), .ZN(n450) );
  XNOR2_X1 U336 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n451) );
  XNOR2_X1 U337 ( .A(n452), .B(n451), .ZN(G1331GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n294) );
  XNOR2_X1 U339 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U341 ( .A(G141GAT), .B(n295), .ZN(n358) );
  XOR2_X1 U342 ( .A(G211GAT), .B(KEYINPUT22), .Z(n297) );
  XNOR2_X1 U343 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT24), .B(KEYINPUT83), .Z(n299) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(G197GAT), .B(KEYINPUT21), .Z(n330) );
  XOR2_X1 U349 ( .A(n300), .B(n330), .Z(n306) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n389) );
  XNOR2_X1 U351 ( .A(G78GAT), .B(G204GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n301), .B(G148GAT), .ZN(n447) );
  XOR2_X1 U353 ( .A(n389), .B(n447), .Z(n303) );
  NAND2_X1 U354 ( .A1(G228GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U356 ( .A(G22GAT), .B(G155GAT), .Z(n407) );
  XNOR2_X1 U357 ( .A(n304), .B(n407), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U359 ( .A(n308), .B(n307), .Z(n309) );
  XNOR2_X1 U360 ( .A(n358), .B(n309), .ZN(n550) );
  XOR2_X1 U361 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(n312), .ZN(n340) );
  XOR2_X1 U365 ( .A(KEYINPUT81), .B(G71GAT), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT80), .B(G176GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n324) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G127GAT), .Z(n408) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G134GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n291), .B(n315), .ZN(n316) );
  NAND2_X1 U371 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n292), .B(n317), .ZN(n318) );
  XOR2_X1 U373 ( .A(n318), .B(G183GAT), .Z(n322) );
  XOR2_X1 U374 ( .A(G120GAT), .B(KEYINPUT79), .Z(n320) );
  XNOR2_X1 U375 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n366) );
  XNOR2_X1 U377 ( .A(n366), .B(KEYINPUT20), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U380 ( .A(n340), .B(n325), .ZN(n555) );
  INV_X1 U381 ( .A(n555), .ZN(n518) );
  XNOR2_X1 U382 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n329), .B(G211GAT), .ZN(n404) );
  XOR2_X1 U386 ( .A(n330), .B(n404), .Z(n332) );
  NAND2_X1 U387 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U389 ( .A(n333), .B(KEYINPUT94), .Z(n336) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n334), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U392 ( .A(n381), .B(KEYINPUT93), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U394 ( .A(G176GAT), .B(G64GAT), .Z(n441) );
  XOR2_X1 U395 ( .A(n337), .B(n441), .Z(n339) );
  XNOR2_X1 U396 ( .A(G204GAT), .B(G92GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n545) );
  XOR2_X1 U399 ( .A(n545), .B(KEYINPUT27), .Z(n373) );
  NAND2_X1 U400 ( .A1(n571), .A2(n373), .ZN(n346) );
  INV_X1 U401 ( .A(n545), .ZN(n483) );
  NAND2_X1 U402 ( .A1(n518), .A2(n483), .ZN(n342) );
  NAND2_X1 U403 ( .A1(n342), .A2(n550), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n343), .B(KEYINPUT25), .ZN(n344) );
  XOR2_X1 U405 ( .A(KEYINPUT98), .B(n344), .Z(n345) );
  NAND2_X1 U406 ( .A1(n346), .A2(n345), .ZN(n371) );
  XOR2_X1 U407 ( .A(G134GAT), .B(KEYINPUT73), .Z(n380) );
  XOR2_X1 U408 ( .A(G85GAT), .B(G155GAT), .Z(n348) );
  XNOR2_X1 U409 ( .A(G29GAT), .B(G162GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U411 ( .A(n380), .B(n349), .Z(n351) );
  NAND2_X1 U412 ( .A1(G225GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n370) );
  XOR2_X1 U414 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n353) );
  XNOR2_X1 U415 ( .A(KEYINPUT92), .B(KEYINPUT88), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U417 ( .A(G57GAT), .B(G148GAT), .Z(n355) );
  XNOR2_X1 U418 ( .A(G1GAT), .B(G127GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U420 ( .A(n357), .B(n356), .Z(n364) );
  INV_X1 U421 ( .A(n358), .ZN(n362) );
  XOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n360) );
  XNOR2_X1 U423 ( .A(KEYINPUT87), .B(KEYINPUT5), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U427 ( .A(n365), .B(KEYINPUT6), .Z(n368) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT1), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U430 ( .A(n370), .B(n369), .Z(n480) );
  INV_X1 U431 ( .A(n480), .ZN(n569) );
  NAND2_X1 U432 ( .A1(n371), .A2(n569), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n372), .B(KEYINPUT99), .ZN(n376) );
  XOR2_X1 U434 ( .A(n550), .B(KEYINPUT28), .Z(n487) );
  NAND2_X1 U435 ( .A1(n480), .A2(n373), .ZN(n533) );
  NOR2_X1 U436 ( .A1(n487), .A2(n533), .ZN(n519) );
  XNOR2_X1 U437 ( .A(n519), .B(KEYINPUT95), .ZN(n374) );
  NOR2_X1 U438 ( .A1(n518), .A2(n374), .ZN(n375) );
  NOR2_X1 U439 ( .A1(n376), .A2(n375), .ZN(n456) );
  XOR2_X1 U440 ( .A(KEYINPUT36), .B(KEYINPUT104), .Z(n400) );
  XOR2_X1 U441 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n378) );
  XNOR2_X1 U442 ( .A(G43GAT), .B(G29GAT), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U444 ( .A(KEYINPUT8), .B(n379), .ZN(n437) );
  INV_X1 U445 ( .A(n437), .ZN(n385) );
  XOR2_X1 U446 ( .A(n381), .B(n380), .Z(n383) );
  NAND2_X1 U447 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT74), .B(KEYINPUT71), .Z(n387) );
  XNOR2_X1 U451 ( .A(KEYINPUT64), .B(KEYINPUT10), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U453 ( .A(n388), .B(KEYINPUT9), .Z(n391) );
  XNOR2_X1 U454 ( .A(n389), .B(KEYINPUT72), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n393) );
  INV_X1 U456 ( .A(KEYINPUT11), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U458 ( .A(G85GAT), .B(G92GAT), .Z(n395) );
  XNOR2_X1 U459 ( .A(G99GAT), .B(G106GAT), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n444) );
  XNOR2_X1 U461 ( .A(n444), .B(KEYINPUT70), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n541) );
  XOR2_X1 U464 ( .A(KEYINPUT75), .B(n541), .Z(n565) );
  XNOR2_X1 U465 ( .A(n400), .B(n565), .ZN(n585) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  INV_X1 U467 ( .A(KEYINPUT14), .ZN(n401) );
  XNOR2_X1 U468 ( .A(G71GAT), .B(G57GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n405), .B(KEYINPUT13), .ZN(n446) );
  XOR2_X1 U470 ( .A(n406), .B(n446), .Z(n410) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U473 ( .A(n411), .B(G64GAT), .Z(n417) );
  XOR2_X1 U474 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n413) );
  XNOR2_X1 U475 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n412) );
  XOR2_X1 U476 ( .A(n413), .B(n412), .Z(n415) );
  XOR2_X1 U477 ( .A(KEYINPUT68), .B(G1GAT), .Z(n431) );
  XNOR2_X1 U478 ( .A(n431), .B(G78GAT), .ZN(n414) );
  INV_X1 U479 ( .A(n581), .ZN(n510) );
  OR2_X1 U480 ( .A1(n456), .A2(n418), .ZN(n419) );
  XNOR2_X1 U481 ( .A(KEYINPUT37), .B(n419), .ZN(n492) );
  XOR2_X1 U482 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n421) );
  XNOR2_X1 U483 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n435) );
  XOR2_X1 U485 ( .A(G22GAT), .B(G141GAT), .Z(n423) );
  XNOR2_X1 U486 ( .A(G50GAT), .B(G36GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U488 ( .A(G113GAT), .B(G15GAT), .Z(n425) );
  XNOR2_X1 U489 ( .A(G169GAT), .B(G197GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U491 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U492 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n429) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U497 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n573) );
  XOR2_X1 U499 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n439) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n578) );
  AND2_X1 U508 ( .A1(n573), .A2(n578), .ZN(n457) );
  XNOR2_X1 U509 ( .A(KEYINPUT38), .B(n450), .ZN(n475) );
  NAND2_X1 U510 ( .A1(n475), .A2(n487), .ZN(n452) );
  OR2_X1 U511 ( .A1(n565), .A2(n510), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n453), .B(KEYINPUT16), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n454), .B(KEYINPUT78), .ZN(n455) );
  NOR2_X1 U514 ( .A1(n456), .A2(n455), .ZN(n478) );
  NAND2_X1 U515 ( .A1(n457), .A2(n478), .ZN(n465) );
  NOR2_X1 U516 ( .A1(n569), .A2(n465), .ZN(n459) );
  XNOR2_X1 U517 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U519 ( .A(G1GAT), .B(n460), .Z(G1324GAT) );
  NOR2_X1 U520 ( .A1(n545), .A2(n465), .ZN(n461) );
  XOR2_X1 U521 ( .A(G8GAT), .B(n461), .Z(G1325GAT) );
  NOR2_X1 U522 ( .A1(n555), .A2(n465), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U525 ( .A(G15GAT), .B(n464), .Z(G1326GAT) );
  INV_X1 U526 ( .A(n487), .ZN(n500) );
  NOR2_X1 U527 ( .A1(n500), .A2(n465), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT102), .B(n466), .Z(n467) );
  XNOR2_X1 U529 ( .A(G22GAT), .B(n467), .ZN(G1327GAT) );
  NAND2_X1 U530 ( .A1(n475), .A2(n480), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n469) );
  XNOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U534 ( .A(KEYINPUT103), .B(n470), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  XOR2_X1 U536 ( .A(G36GAT), .B(KEYINPUT107), .Z(n474) );
  NAND2_X1 U537 ( .A1(n475), .A2(n483), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n474), .B(n473), .ZN(G1329GAT) );
  NAND2_X1 U539 ( .A1(n475), .A2(n518), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n476), .B(KEYINPUT40), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n477), .B(G43GAT), .ZN(G1330GAT) );
  XNOR2_X1 U542 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n482) );
  XOR2_X1 U543 ( .A(n578), .B(KEYINPUT41), .Z(n503) );
  NOR2_X1 U544 ( .A1(n573), .A2(n503), .ZN(n491) );
  NAND2_X1 U545 ( .A1(n478), .A2(n491), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n479), .B(KEYINPUT109), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n480), .A2(n488), .ZN(n481) );
  XNOR2_X1 U548 ( .A(n482), .B(n481), .ZN(G1332GAT) );
  NAND2_X1 U549 ( .A1(n483), .A2(n488), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n484), .B(KEYINPUT110), .ZN(n485) );
  XNOR2_X1 U551 ( .A(G64GAT), .B(n485), .ZN(G1333GAT) );
  NAND2_X1 U552 ( .A1(n518), .A2(n488), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n486), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U554 ( .A(G78GAT), .B(KEYINPUT43), .Z(n490) );
  NAND2_X1 U555 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n490), .B(n489), .ZN(G1335GAT) );
  NAND2_X1 U557 ( .A1(n492), .A2(n491), .ZN(n499) );
  NOR2_X1 U558 ( .A1(n569), .A2(n499), .ZN(n494) );
  XNOR2_X1 U559 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n493) );
  XNOR2_X1 U560 ( .A(n494), .B(n493), .ZN(G1336GAT) );
  NOR2_X1 U561 ( .A1(n545), .A2(n499), .ZN(n495) );
  XOR2_X1 U562 ( .A(G92GAT), .B(n495), .Z(G1337GAT) );
  NOR2_X1 U563 ( .A1(n555), .A2(n499), .ZN(n496) );
  XOR2_X1 U564 ( .A(G99GAT), .B(n496), .Z(G1338GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n498) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n497) );
  XNOR2_X1 U567 ( .A(n498), .B(n497), .ZN(n502) );
  NOR2_X1 U568 ( .A1(n500), .A2(n499), .ZN(n501) );
  XOR2_X1 U569 ( .A(n502), .B(n501), .Z(G1339GAT) );
  XNOR2_X1 U570 ( .A(n581), .B(KEYINPUT114), .ZN(n562) );
  XOR2_X1 U571 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n505) );
  INV_X1 U572 ( .A(n503), .ZN(n557) );
  NAND2_X1 U573 ( .A1(n557), .A2(n573), .ZN(n504) );
  XOR2_X1 U574 ( .A(n505), .B(n504), .Z(n506) );
  OR2_X1 U575 ( .A1(n562), .A2(n506), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n507), .B(KEYINPUT116), .ZN(n508) );
  NOR2_X1 U577 ( .A1(n541), .A2(n508), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n509), .B(KEYINPUT47), .ZN(n516) );
  NOR2_X1 U579 ( .A1(n585), .A2(n510), .ZN(n511) );
  XNOR2_X1 U580 ( .A(KEYINPUT45), .B(n511), .ZN(n512) );
  NAND2_X1 U581 ( .A1(n512), .A2(n578), .ZN(n513) );
  NOR2_X1 U582 ( .A1(n573), .A2(n513), .ZN(n514) );
  XNOR2_X1 U583 ( .A(KEYINPUT117), .B(n514), .ZN(n515) );
  AND2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(KEYINPUT48), .ZN(n546) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U587 ( .A1(n546), .A2(n520), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n527), .A2(n573), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n523) );
  NAND2_X1 U591 ( .A1(n527), .A2(n557), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n524), .ZN(G1341GAT) );
  NAND2_X1 U594 ( .A1(n562), .A2(n527), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n525), .B(KEYINPUT50), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n526), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n529) );
  NAND2_X1 U598 ( .A1(n527), .A2(n565), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U600 ( .A(G134GAT), .B(n530), .Z(G1343GAT) );
  INV_X1 U601 ( .A(n546), .ZN(n531) );
  NAND2_X1 U602 ( .A1(n531), .A2(n571), .ZN(n532) );
  NOR2_X1 U603 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n573), .A2(n542), .ZN(n534) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n534), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n536) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n535) );
  XNOR2_X1 U608 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(n537), .Z(n539) );
  NAND2_X1 U610 ( .A1(n542), .A2(n557), .ZN(n538) );
  XNOR2_X1 U611 ( .A(n539), .B(n538), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n542), .A2(n581), .ZN(n540) );
  XNOR2_X1 U613 ( .A(n540), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U615 ( .A(n543), .B(KEYINPUT122), .ZN(n544) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n544), .ZN(G1347GAT) );
  NOR2_X1 U617 ( .A1(n546), .A2(n545), .ZN(n549) );
  INV_X1 U618 ( .A(KEYINPUT54), .ZN(n547) );
  AND2_X1 U619 ( .A1(n569), .A2(n550), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n570), .A2(n551), .ZN(n553) );
  XOR2_X1 U621 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n566), .A2(n573), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n566), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT125), .Z(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n562), .A2(n566), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT126), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .Z(n575) );
  AND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  INV_X1 U639 ( .A(n584), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(KEYINPUT127), .Z(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  OR2_X1 U645 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

