//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n204), .A3(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n197), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n201), .A2(G134), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n199), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G128), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT64), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n192), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G128), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n212), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(new_n208), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n212), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(G143), .B2(new_n188), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n217), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n219), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n222), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n195), .A2(new_n196), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n207), .A2(new_n205), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G119), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT65), .A3(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(G119), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT2), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT2), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G113), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n247), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(new_n239), .A3(new_n241), .A4(new_n242), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT68), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(new_n249), .B2(new_n251), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n221), .A2(new_n236), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n207), .A2(new_n205), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(new_n197), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT66), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(new_n254), .A3(new_n231), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n249), .A2(new_n251), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n208), .B2(new_n220), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT28), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n258), .A2(new_n260), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n216), .A2(new_n219), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(new_n222), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n263), .A2(new_n281), .A3(new_n264), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n279), .B1(new_n208), .B2(new_n220), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n266), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n266), .A4(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n265), .A2(new_n276), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT31), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n292), .B(new_n289), .C1(new_n286), .C2(new_n287), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n278), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G472), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n288), .A2(new_n265), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n277), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n277), .B1(new_n268), .B2(KEYINPUT28), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n258), .A3(new_n260), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n304), .A2(new_n258), .A3(new_n308), .A4(new_n260), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n303), .A2(new_n306), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n260), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n263), .A2(new_n231), .A3(new_n264), .ZN(new_n314));
  INV_X1    g128(.A(new_n254), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n256), .B1(new_n316), .B2(new_n265), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n259), .B1(new_n255), .B2(new_n256), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n313), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n277), .A2(new_n307), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n301), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n187), .B1(new_n300), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT32), .B1(new_n294), .B2(new_n295), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n322), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G217), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n311), .B2(G234), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  OR3_X1    g150(.A1(new_n336), .A2(KEYINPUT16), .A3(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(G146), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n188), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n240), .B2(G128), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n341), .B(new_n342), .C1(G119), .C2(new_n223), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n343), .A2(G110), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  XNOR2_X1  g159(.A(G119), .B(G128), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT24), .B(G110), .Z(new_n347));
  OAI22_X1  g161(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n344), .A2(new_n345), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n338), .B(new_n339), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n346), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n353), .A3(new_n346), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n352), .A2(new_n354), .B1(G110), .B2(new_n343), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n335), .A2(new_n337), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n188), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n338), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n355), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n350), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT77), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G137), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n350), .B(new_n366), .C1(new_n360), .C2(new_n361), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n333), .B1(new_n370), .B2(new_n312), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n368), .A2(KEYINPUT25), .A3(new_n311), .A4(new_n369), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n332), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n331), .A2(G902), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT78), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g191(.A(KEYINPUT84), .B(G469), .Z(new_n378));
  AND2_X1   g192(.A1(new_n234), .A2(KEYINPUT82), .ZN(new_n379));
  INV_X1    g193(.A(G101), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G104), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(KEYINPUT79), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(KEYINPUT80), .A3(G104), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n386), .B2(new_n387), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n380), .B(new_n385), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n384), .B2(new_n382), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n280), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n192), .B1(new_n224), .B2(new_n223), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n219), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n379), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT82), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT12), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  OAI221_X1 g216(.A(new_n379), .B1(KEYINPUT12), .B2(new_n400), .C1(new_n393), .C2(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  INV_X1    g219(.A(G227), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n405), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT81), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(G101), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n233), .B1(new_n413), .B2(KEYINPUT4), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n280), .A2(KEYINPUT10), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n391), .A2(new_n392), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n424), .B1(new_n425), .B2(new_n396), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n262), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n404), .A2(new_n409), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n410), .B1(KEYINPUT81), .B2(new_n413), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n418), .B1(new_n429), .B2(new_n416), .ZN(new_n430));
  OAI22_X1  g244(.A1(new_n397), .A2(KEYINPUT10), .B1(new_n421), .B2(new_n423), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n234), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n409), .B1(new_n432), .B2(new_n427), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n428), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g249(.A(KEYINPUT85), .B(new_n409), .C1(new_n432), .C2(new_n427), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n311), .B(new_n378), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n404), .A2(KEYINPUT83), .A3(new_n427), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT83), .B1(new_n404), .B2(new_n427), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n408), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n427), .A2(new_n409), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n432), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n437), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT9), .B(G234), .ZN(new_n447));
  OAI21_X1  g261(.A(G221), .B1(new_n447), .B2(G902), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n266), .B1(new_n413), .B2(KEYINPUT4), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n429), .B2(new_n416), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(G116), .A3(new_n240), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G113), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n243), .A2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n251), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n423), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n452), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  INV_X1    g276(.A(new_n417), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n462), .B(new_n451), .C1(new_n463), .C2(new_n453), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n464), .A3(KEYINPUT6), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n452), .C1(new_n454), .C2(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n197), .A2(G125), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n216), .A2(new_n336), .A3(new_n219), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n272), .A2(G224), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n472), .B(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT88), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n243), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n251), .B1(new_n457), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n424), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n451), .B(KEYINPUT8), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n483), .B(new_n484), .C1(new_n424), .C2(new_n459), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n470), .A2(new_n468), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n474), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n474), .A2(new_n487), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n491), .B2(new_n464), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n476), .A2(new_n479), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n479), .B1(new_n476), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n450), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n449), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n334), .A2(KEYINPUT90), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n336), .A2(G140), .ZN(new_n500));
  INV_X1    g314(.A(G140), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G125), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n498), .A2(new_n503), .A3(G146), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n339), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n190), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n271), .A2(new_n272), .A3(G143), .A4(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n509), .A2(KEYINPUT89), .A3(new_n510), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT89), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n505), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT19), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT19), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n334), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n498), .A2(new_n503), .A3(new_n516), .A4(KEYINPUT19), .ZN(new_n520));
  AOI21_X1  g334(.A(G146), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n509), .A2(G131), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n507), .A2(new_n203), .A3(new_n508), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n338), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n514), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n383), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n522), .A2(new_n531), .A3(new_n523), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n509), .A2(KEYINPUT17), .A3(G131), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n357), .A3(new_n338), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n514), .A3(new_n528), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n530), .B2(new_n535), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n537), .A2(new_n539), .B1(new_n541), .B2(KEYINPUT20), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n536), .A2(new_n540), .A3(new_n543), .A4(new_n538), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n535), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n528), .B1(new_n534), .B2(new_n514), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G475), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT13), .B1(new_n223), .B2(G143), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n199), .ZN(new_n553));
  XNOR2_X1  g367(.A(G128), .B(G143), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G116), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n238), .A2(G122), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n381), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n381), .B1(new_n559), .B2(new_n560), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n555), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n557), .B(KEYINPUT93), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n560), .B(KEYINPUT14), .ZN(new_n566));
  OAI21_X1  g380(.A(G107), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n554), .B(new_n199), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n561), .A3(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n447), .A2(new_n330), .A3(G953), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n564), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n311), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n573), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n272), .B(new_n311), .C1(G234), .C2(G237), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT21), .B(G898), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G952), .ZN(new_n581));
  AOI211_X1 g395(.A(G953), .B(new_n581), .C1(G234), .C2(G237), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT94), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n551), .A2(new_n577), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n329), .A2(new_n377), .A3(new_n497), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  AND3_X1   g403(.A1(new_n476), .A2(new_n477), .A3(new_n492), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n477), .B1(new_n476), .B2(new_n492), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n450), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR3_X1    g406(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT33), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT33), .B1(new_n571), .B2(new_n572), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n312), .A2(new_n574), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n595), .A2(new_n596), .B1(new_n574), .B2(new_n573), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n551), .A2(new_n585), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT95), .B1(new_n592), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n450), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n476), .A2(new_n492), .ZN(new_n602));
  INV_X1    g416(.A(new_n477), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n476), .A2(new_n477), .A3(new_n492), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n542), .A2(new_n544), .B1(G475), .B2(new_n549), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n608), .A2(new_n586), .A3(new_n597), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n377), .ZN(new_n612));
  INV_X1    g426(.A(new_n296), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n301), .B1(new_n294), .B2(new_n311), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n448), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n404), .A2(new_n427), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n438), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(new_n408), .B1(new_n442), .B2(new_n432), .ZN(new_n621));
  OAI21_X1  g435(.A(G469), .B1(new_n621), .B2(G902), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n616), .B1(new_n622), .B2(new_n437), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n611), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  AOI21_X1  g441(.A(new_n543), .B1(new_n536), .B2(new_n538), .ZN(new_n628));
  AOI211_X1 g442(.A(KEYINPUT20), .B(new_n539), .C1(new_n530), .C2(new_n535), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n550), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n576), .A2(new_n630), .A3(new_n586), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n631), .B(new_n450), .C1(new_n591), .C2(new_n590), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NAND2_X1  g449(.A1(new_n294), .A2(new_n311), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n371), .A2(new_n372), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n331), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n362), .B(new_n640), .Z(new_n641));
  INV_X1    g455(.A(new_n375), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n637), .A2(new_n587), .A3(new_n644), .A4(new_n296), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n645), .A2(new_n449), .A3(new_n496), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  NAND3_X1  g462(.A1(new_n446), .A2(new_n448), .A3(new_n644), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n323), .B2(new_n328), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n578), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n583), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n576), .A2(new_n630), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n606), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XNOR2_X1  g473(.A(new_n653), .B(KEYINPUT39), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n623), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT98), .Z(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n664));
  INV_X1    g478(.A(new_n316), .ZN(new_n665));
  INV_X1    g479(.A(new_n265), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n546), .B1(new_n668), .B2(new_n276), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n277), .B1(new_n288), .B2(new_n265), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n326), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT97), .Z(new_n673));
  INV_X1    g487(.A(new_n495), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n493), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n608), .A2(new_n576), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n644), .A2(new_n601), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n663), .A2(new_n664), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  INV_X1    g497(.A(new_n649), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n551), .A2(new_n598), .A3(new_n653), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n592), .A2(new_n685), .A3(KEYINPUT99), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n608), .A2(new_n597), .A3(new_n654), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n606), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n329), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n650), .A2(KEYINPUT100), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT101), .B(G146), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G48));
  NOR3_X1   g511(.A1(new_n430), .A2(new_n234), .A3(new_n431), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n262), .B1(new_n420), .B2(new_n426), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n408), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n700), .A2(KEYINPUT85), .B1(new_n442), .B2(new_n404), .ZN(new_n701));
  INV_X1    g515(.A(new_n436), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n312), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n448), .B(new_n437), .C1(new_n703), .C2(new_n445), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n311), .B1(new_n435), .B2(new_n436), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n448), .A4(new_n437), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n600), .A2(new_n610), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n329), .A2(new_n711), .A3(new_n377), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  INV_X1    g529(.A(new_n632), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n705), .A2(new_n716), .A3(new_n709), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n329), .A2(new_n717), .A3(new_n377), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  OR2_X1    g533(.A1(new_n704), .A2(new_n592), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n587), .A2(new_n644), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n329), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND2_X1  g538(.A1(new_n606), .A2(new_n678), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n705), .A3(new_n585), .A4(new_n709), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI22_X1  g542(.A1(new_n291), .A2(new_n293), .B1(new_n319), .B2(new_n276), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n295), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(KEYINPUT103), .A3(new_n295), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n614), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n614), .A2(new_n734), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n376), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT105), .B1(new_n639), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n373), .A2(new_n741), .A3(new_n376), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT106), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n740), .A2(new_n742), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n735), .A2(new_n745), .A3(new_n737), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n728), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  INV_X1    g563(.A(new_n733), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT103), .B1(new_n729), .B2(new_n295), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n637), .A2(KEYINPUT104), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n644), .A4(new_n736), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n707), .A2(new_n437), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n448), .A3(new_n606), .A4(new_n688), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n336), .ZN(G27));
  OR2_X1    g572(.A1(new_n299), .A2(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n299), .A2(KEYINPUT107), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n327), .A3(new_n298), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n743), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n674), .A2(new_n450), .A3(new_n493), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n623), .A2(KEYINPUT42), .A3(new_n688), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n449), .A2(new_n763), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n329), .A2(new_n377), .A3(new_n688), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n203), .ZN(G33));
  AOI21_X1  g585(.A(new_n612), .B1(new_n323), .B2(new_n328), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n655), .A3(new_n767), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NAND2_X1  g588(.A1(new_n441), .A2(new_n443), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n445), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  NAND2_X1  g592(.A1(G469), .A2(G902), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n779), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n437), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n448), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n660), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n598), .A2(new_n608), .ZN(new_n788));
  NAND2_X1  g602(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n644), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n613), .A2(new_n614), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n764), .A3(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  OAI21_X1  g614(.A(new_n785), .B1(KEYINPUT109), .B2(KEYINPUT47), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n329), .A2(new_n377), .A3(new_n685), .A4(new_n763), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n803));
  OAI211_X1 g617(.A(new_n801), .B(new_n802), .C1(new_n785), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT110), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NOR4_X1   g620(.A1(new_n745), .A2(new_n601), .A3(new_n616), .A4(new_n788), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n755), .B(KEYINPUT49), .ZN(new_n808));
  INV_X1    g622(.A(new_n677), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n673), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n757), .B1(new_n650), .B2(new_n657), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n653), .B(KEYINPUT114), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n449), .A2(new_n644), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n672), .A3(new_n726), .ZN(new_n814));
  AND4_X1   g628(.A1(KEYINPUT100), .A2(new_n329), .A3(new_n684), .A4(new_n690), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT100), .B1(new_n650), .B2(new_n690), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n811), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n695), .A2(KEYINPUT52), .A3(new_n811), .A4(new_n814), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n713), .A2(new_n718), .A3(new_n723), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n743), .A2(new_n736), .A3(new_n753), .A4(new_n752), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n746), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n738), .A2(KEYINPUT106), .A3(new_n743), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n727), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n770), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n738), .A2(new_n767), .A3(new_n644), .A4(new_n688), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n763), .A2(new_n577), .A3(new_n630), .A4(new_n654), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n329), .A2(new_n684), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n773), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n601), .B1(new_n674), .B2(new_n493), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n446), .A2(new_n834), .A3(new_n448), .A4(new_n587), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n612), .B(new_n835), .C1(new_n323), .C2(new_n328), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n637), .A2(new_n296), .A3(new_n377), .A4(new_n609), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n645), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n497), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n551), .A2(new_n576), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n585), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT111), .B1(new_n841), .B2(new_n496), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n834), .A2(new_n843), .A3(new_n585), .A4(new_n840), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n615), .A3(new_n844), .A4(new_n623), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT112), .B1(new_n836), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n588), .A2(new_n848), .A3(new_n839), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n773), .A2(KEYINPUT113), .A3(new_n828), .A4(new_n830), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n827), .A2(new_n833), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n821), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n833), .A3(new_n851), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n822), .A2(new_n826), .ZN(new_n856));
  INV_X1    g670(.A(new_n770), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n819), .A2(new_n820), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n853), .B1(new_n821), .B2(new_n852), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  AND4_X1   g678(.A1(KEYINPUT53), .A2(new_n850), .A3(new_n833), .A4(new_n851), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n611), .A2(new_n710), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n867), .A2(new_n772), .B1(new_n329), .B2(new_n722), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n748), .A2(new_n868), .A3(new_n718), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n869), .B2(new_n770), .ZN(new_n870));
  INV_X1    g684(.A(new_n822), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n857), .A2(new_n871), .A3(KEYINPUT115), .A4(new_n748), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n865), .A2(new_n860), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n864), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n704), .A2(new_n763), .A3(new_n583), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n792), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT118), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n644), .A3(new_n738), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n876), .A2(new_n377), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n673), .A2(new_n608), .A3(new_n597), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n755), .A2(new_n616), .ZN(new_n883));
  INV_X1    g697(.A(new_n801), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n785), .A2(new_n803), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n824), .A2(new_n825), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n792), .A2(new_n582), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n763), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n882), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n677), .A2(new_n450), .A3(new_n704), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT50), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n894), .B(new_n896), .Z(new_n897));
  AOI21_X1  g711(.A(KEYINPUT116), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n581), .A2(G953), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n608), .A2(new_n597), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n673), .A2(new_n902), .A3(new_n880), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n901), .B(new_n903), .C1(new_n890), .C2(new_n720), .ZN(new_n904));
  INV_X1    g718(.A(new_n762), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n878), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT48), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n906), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(KEYINPUT48), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n898), .B2(new_n899), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n875), .A2(new_n900), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n810), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NAND2_X1  g729(.A1(new_n863), .A2(new_n873), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n312), .A3(new_n603), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n465), .A2(new_n467), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n475), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT55), .Z(new_n920));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(KEYINPUT56), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n272), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  XOR2_X1   g740(.A(new_n779), .B(KEYINPUT57), .Z(new_n927));
  INV_X1    g741(.A(new_n874), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n864), .B1(new_n863), .B2(new_n873), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n436), .B2(new_n435), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n916), .A2(new_n312), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(new_n778), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n925), .B1(new_n931), .B2(new_n933), .ZN(G54));
  NAND2_X1  g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT121), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n537), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n925), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n916), .A2(new_n312), .A3(new_n536), .A4(new_n936), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT59), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n595), .B(new_n944), .C1(new_n928), .C2(new_n929), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n939), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n595), .B1(new_n875), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n870), .A2(new_n872), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n850), .A2(new_n833), .A3(KEYINPUT53), .A4(new_n851), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n821), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(new_n861), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n925), .B1(new_n955), .B2(new_n370), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n957));
  AND4_X1   g771(.A1(new_n957), .A2(new_n916), .A3(new_n641), .A4(new_n951), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n950), .B1(new_n863), .B2(new_n873), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(new_n641), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n956), .B(KEYINPUT61), .C1(new_n958), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  INV_X1    g779(.A(new_n579), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n272), .B1(new_n966), .B2(G224), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n850), .A2(new_n856), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT123), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n272), .ZN(new_n970));
  INV_X1    g784(.A(G898), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n918), .B1(new_n971), .B2(G953), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  OAI21_X1  g787(.A(G953), .B1(new_n406), .B2(new_n651), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n282), .A2(new_n283), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n519), .A2(new_n520), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n974), .B1(new_n978), .B2(KEYINPUT125), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n660), .A2(new_n786), .A3(new_n726), .A4(new_n905), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT124), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n695), .A2(new_n811), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n799), .A2(new_n857), .A3(new_n773), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n805), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n985), .A2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n978), .B1(new_n651), .B2(new_n272), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n682), .A2(new_n983), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n772), .B(new_n764), .C1(new_n902), .C2(new_n840), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n662), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n799), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(new_n805), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n272), .ZN(new_n995));
  OAI221_X1 g809(.A(new_n980), .B1(new_n986), .B2(new_n987), .C1(new_n995), .C2(new_n978), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n986), .A2(new_n987), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n978), .B1(new_n994), .B2(new_n272), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n979), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(new_n999), .ZN(G72));
  XNOR2_X1  g814(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n301), .A2(new_n546), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n994), .B2(new_n969), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n925), .B1(new_n1005), .B2(new_n670), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n288), .A2(new_n290), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n303), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n854), .B2(new_n861), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1004), .B1(new_n985), .B2(new_n969), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1010), .A2(new_n277), .A3(new_n265), .A4(new_n288), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1006), .A2(new_n1009), .A3(new_n1011), .ZN(G57));
endmodule


