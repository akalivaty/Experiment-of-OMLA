

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n555), .A2(n524), .ZN(n763) );
  XOR2_X1 U553 ( .A(KEYINPUT15), .B(n658), .Z(n944) );
  XNOR2_X1 U554 ( .A(KEYINPUT30), .B(KEYINPUT92), .ZN(n678) );
  NAND2_X1 U555 ( .A1(n660), .A2(n659), .ZN(n661) );
  INV_X1 U556 ( .A(n944), .ZN(n659) );
  INV_X1 U557 ( .A(KEYINPUT32), .ZN(n537) );
  NAND2_X1 U558 ( .A1(n519), .A2(n528), .ZN(n724) );
  NAND2_X1 U559 ( .A1(n531), .A2(n529), .ZN(n528) );
  NOR2_X1 U560 ( .A1(n701), .A2(n549), .ZN(n545) );
  AND2_X1 U561 ( .A1(n748), .A2(n746), .ZN(n672) );
  NAND2_X1 U562 ( .A1(n554), .A2(n664), .ZN(n553) );
  NOR2_X1 U563 ( .A1(n669), .A2(n518), .ZN(n554) );
  AND2_X1 U564 ( .A1(n648), .A2(n647), .ZN(n662) );
  XNOR2_X1 U565 ( .A(n551), .B(n550), .ZN(n676) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n550) );
  NAND2_X1 U567 ( .A1(n553), .A2(n552), .ZN(n551) );
  XNOR2_X1 U568 ( .A(n671), .B(KEYINPUT28), .ZN(n552) );
  AND2_X1 U569 ( .A1(n677), .A2(n547), .ZN(n701) );
  AND2_X1 U570 ( .A1(n548), .A2(G8), .ZN(n547) );
  INV_X1 U571 ( .A(G1966), .ZN(n548) );
  NAND2_X1 U572 ( .A1(n537), .A2(n549), .ZN(n536) );
  AND2_X1 U573 ( .A1(n530), .A2(KEYINPUT97), .ZN(n529) );
  AND2_X1 U574 ( .A1(n725), .A2(n691), .ZN(n726) );
  XNOR2_X1 U575 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n627) );
  INV_X1 U576 ( .A(n627), .ZN(n544) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n748) );
  NOR2_X1 U578 ( .A1(n606), .A2(n565), .ZN(n810) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n566), .Z(n811) );
  AND2_X1 U580 ( .A1(G2104), .A2(n578), .ZN(n575) );
  NOR2_X2 U581 ( .A1(G2104), .A2(n578), .ZN(n898) );
  NAND2_X1 U582 ( .A1(n544), .A2(n543), .ZN(n542) );
  INV_X1 U583 ( .A(G101), .ZN(n543) );
  NOR2_X1 U584 ( .A1(n763), .A2(n762), .ZN(n765) );
  NOR2_X1 U585 ( .A1(n606), .A2(G651), .ZN(n818) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n814) );
  XNOR2_X1 U587 ( .A(n574), .B(n573), .ZN(n901) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n574) );
  XNOR2_X1 U589 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U590 ( .A1(n677), .A2(G8), .ZN(n691) );
  AND2_X1 U591 ( .A1(n663), .A2(n944), .ZN(n518) );
  AND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n519) );
  NOR2_X1 U593 ( .A1(n782), .A2(n632), .ZN(n520) );
  AND2_X1 U594 ( .A1(n704), .A2(n536), .ZN(n521) );
  AND2_X1 U595 ( .A1(n628), .A2(n542), .ZN(n522) );
  NAND2_X1 U596 ( .A1(n627), .A2(G101), .ZN(n523) );
  OR2_X1 U597 ( .A1(n691), .A2(n728), .ZN(n524) );
  AND2_X1 U598 ( .A1(n633), .A2(n520), .ZN(n746) );
  AND2_X1 U599 ( .A1(n537), .A2(n705), .ZN(n525) );
  AND2_X1 U600 ( .A1(KEYINPUT32), .A2(G8), .ZN(n526) );
  INV_X1 U601 ( .A(n687), .ZN(n700) );
  NAND2_X1 U602 ( .A1(n699), .A2(n527), .ZN(n687) );
  XNOR2_X1 U603 ( .A(n686), .B(KEYINPUT31), .ZN(n527) );
  NAND2_X1 U604 ( .A1(n534), .A2(n537), .ZN(n530) );
  INV_X1 U605 ( .A(n535), .ZN(n531) );
  NAND2_X1 U606 ( .A1(n534), .A2(n525), .ZN(n532) );
  NAND2_X1 U607 ( .A1(n535), .A2(n705), .ZN(n533) );
  INV_X1 U608 ( .A(n697), .ZN(n534) );
  NAND2_X1 U609 ( .A1(n538), .A2(n521), .ZN(n535) );
  NAND2_X1 U610 ( .A1(n697), .A2(n526), .ZN(n538) );
  NAND2_X1 U611 ( .A1(n522), .A2(n539), .ZN(n629) );
  NAND2_X1 U612 ( .A1(n541), .A2(n540), .ZN(n539) );
  NAND2_X1 U613 ( .A1(n902), .A2(n523), .ZN(n540) );
  OR2_X1 U614 ( .A1(n902), .A2(n544), .ZN(n541) );
  XNOR2_X2 U615 ( .A(n575), .B(KEYINPUT64), .ZN(n902) );
  INV_X1 U616 ( .A(n698), .ZN(n546) );
  NAND2_X1 U617 ( .A1(n546), .A2(n545), .ZN(n679) );
  INV_X1 U618 ( .A(G8), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT103), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n559), .A2(n557), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n726), .B(n558), .ZN(n557) );
  INV_X1 U622 ( .A(KEYINPUT102), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n720), .A2(n719), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n672), .A2(G2072), .ZN(n666) );
  AND2_X1 U625 ( .A1(n672), .A2(G1996), .ZN(n634) );
  INV_X1 U626 ( .A(KEYINPUT27), .ZN(n665) );
  XNOR2_X1 U627 ( .A(n666), .B(n665), .ZN(n668) );
  INV_X1 U628 ( .A(KEYINPUT95), .ZN(n688) );
  INV_X1 U629 ( .A(KEYINPUT97), .ZN(n705) );
  INV_X1 U630 ( .A(G40), .ZN(n632) );
  INV_X1 U631 ( .A(n746), .ZN(n747) );
  INV_X1 U632 ( .A(G2105), .ZN(n578) );
  INV_X1 U633 ( .A(KEYINPUT17), .ZN(n573) );
  INV_X1 U634 ( .A(KEYINPUT104), .ZN(n764) );
  XNOR2_X1 U635 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n780) );
  XOR2_X1 U636 ( .A(KEYINPUT0), .B(G543), .Z(n606) );
  INV_X1 U637 ( .A(G651), .ZN(n565) );
  NAND2_X1 U638 ( .A1(n810), .A2(G76), .ZN(n560) );
  XNOR2_X1 U639 ( .A(KEYINPUT72), .B(n560), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n814), .A2(G89), .ZN(n561) );
  XNOR2_X1 U641 ( .A(KEYINPUT4), .B(n561), .ZN(n562) );
  NAND2_X1 U642 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U643 ( .A(n564), .B(KEYINPUT5), .ZN(n571) );
  NOR2_X1 U644 ( .A1(G543), .A2(n565), .ZN(n566) );
  NAND2_X1 U645 ( .A1(G63), .A2(n811), .ZN(n568) );
  NAND2_X1 U646 ( .A1(G51), .A2(n818), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U648 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U649 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U650 ( .A1(G138), .A2(n901), .ZN(n577) );
  NAND2_X1 U651 ( .A1(G102), .A2(n902), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n582) );
  AND2_X1 U653 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U654 ( .A1(G114), .A2(n897), .ZN(n580) );
  NAND2_X1 U655 ( .A1(G126), .A2(n898), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U657 ( .A1(n582), .A2(n581), .ZN(G164) );
  NAND2_X1 U658 ( .A1(G65), .A2(n811), .ZN(n584) );
  NAND2_X1 U659 ( .A1(G53), .A2(n818), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT68), .B(n585), .Z(n589) );
  NAND2_X1 U662 ( .A1(G91), .A2(n814), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G78), .A2(n810), .ZN(n586) );
  AND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(G299) );
  NAND2_X1 U666 ( .A1(G64), .A2(n811), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G52), .A2(n818), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U669 ( .A(KEYINPUT67), .B(n592), .Z(n597) );
  NAND2_X1 U670 ( .A1(G90), .A2(n814), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G77), .A2(n810), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U673 ( .A(KEYINPUT9), .B(n595), .Z(n596) );
  NOR2_X1 U674 ( .A1(n597), .A2(n596), .ZN(G171) );
  INV_X1 U675 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U676 ( .A(G168), .B(KEYINPUT8), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n598), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U678 ( .A1(G88), .A2(n814), .ZN(n600) );
  NAND2_X1 U679 ( .A1(G75), .A2(n810), .ZN(n599) );
  NAND2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U681 ( .A(KEYINPUT81), .B(n601), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G62), .A2(n811), .ZN(n603) );
  NAND2_X1 U683 ( .A1(G50), .A2(n818), .ZN(n602) );
  AND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(G303) );
  NAND2_X1 U686 ( .A1(G87), .A2(n606), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G49), .A2(n818), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G74), .A2(G651), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U690 ( .A1(n811), .A2(n609), .ZN(n610) );
  XOR2_X1 U691 ( .A(KEYINPUT79), .B(n610), .Z(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(n613), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U694 ( .A1(G86), .A2(n814), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G61), .A2(n811), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n810), .A2(G73), .ZN(n616) );
  XOR2_X1 U698 ( .A(KEYINPUT2), .B(n616), .Z(n617) );
  NOR2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n818), .A2(G48), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(G305) );
  INV_X1 U702 ( .A(G303), .ZN(G166) );
  NAND2_X1 U703 ( .A1(G85), .A2(n814), .ZN(n622) );
  NAND2_X1 U704 ( .A1(G72), .A2(n810), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G60), .A2(n811), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G47), .A2(n818), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(G290) );
  NAND2_X1 U710 ( .A1(G125), .A2(n898), .ZN(n628) );
  XNOR2_X1 U711 ( .A(n629), .B(KEYINPUT66), .ZN(n783) );
  INV_X1 U712 ( .A(n783), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G137), .A2(n901), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G113), .A2(n897), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n782) );
  XOR2_X1 U716 ( .A(n634), .B(KEYINPUT26), .Z(n648) );
  NAND2_X2 U717 ( .A1(n748), .A2(n746), .ZN(n677) );
  NAND2_X1 U718 ( .A1(n677), .A2(G1341), .ZN(n646) );
  NAND2_X1 U719 ( .A1(G68), .A2(n810), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n814), .A2(G81), .ZN(n635) );
  XNOR2_X1 U721 ( .A(n635), .B(KEYINPUT12), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n638) );
  XNOR2_X1 U724 ( .A(n639), .B(n638), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n811), .A2(G56), .ZN(n640) );
  XOR2_X1 U726 ( .A(KEYINPUT14), .B(n640), .Z(n641) );
  NOR2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n818), .A2(G43), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n941) );
  INV_X1 U730 ( .A(n941), .ZN(n645) );
  AND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G1348), .A2(n677), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n672), .A2(G2067), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U735 ( .A(KEYINPUT91), .B(n651), .ZN(n663) );
  INV_X1 U736 ( .A(n663), .ZN(n660) );
  NAND2_X1 U737 ( .A1(G92), .A2(n814), .ZN(n653) );
  NAND2_X1 U738 ( .A1(G79), .A2(n810), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U740 ( .A1(G66), .A2(n811), .ZN(n655) );
  NAND2_X1 U741 ( .A1(G54), .A2(n818), .ZN(n654) );
  NAND2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U744 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G1956), .A2(n677), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n670) );
  NOR2_X1 U747 ( .A1(n670), .A2(G299), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G299), .A2(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G1961), .A2(n677), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT25), .B(G2078), .Z(n1026) );
  NAND2_X1 U751 ( .A1(n672), .A2(n1026), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n682) );
  OR2_X1 U753 ( .A1(n682), .A2(G301), .ZN(n675) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n699) );
  NOR2_X1 U755 ( .A1(G2084), .A2(n677), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n680), .A2(G168), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(KEYINPUT93), .ZN(n685) );
  NAND2_X1 U759 ( .A1(G301), .A2(n682), .ZN(n683) );
  XNOR2_X1 U760 ( .A(KEYINPUT94), .B(n683), .ZN(n684) );
  NAND2_X1 U761 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U762 ( .A1(n687), .A2(G286), .ZN(n689) );
  XNOR2_X1 U763 ( .A(n689), .B(n688), .ZN(n696) );
  NOR2_X1 U764 ( .A1(G2090), .A2(n677), .ZN(n690) );
  XNOR2_X1 U765 ( .A(n690), .B(KEYINPUT96), .ZN(n693) );
  NOR2_X1 U766 ( .A1(n691), .A2(G1971), .ZN(n692) );
  NOR2_X1 U767 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U768 ( .A1(G303), .A2(n694), .ZN(n695) );
  NAND2_X1 U769 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U770 ( .A1(G8), .A2(n698), .ZN(n703) );
  NOR2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U773 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NOR2_X1 U774 ( .A1(G1971), .A2(G303), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n706), .B(KEYINPUT98), .ZN(n707) );
  NOR2_X1 U776 ( .A1(n958), .A2(n707), .ZN(n709) );
  INV_X1 U777 ( .A(KEYINPUT33), .ZN(n708) );
  AND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n724), .A2(n710), .ZN(n714) );
  INV_X1 U780 ( .A(n691), .ZN(n711) );
  NAND2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n959) );
  AND2_X1 U782 ( .A1(n711), .A2(n959), .ZN(n712) );
  OR2_X1 U783 ( .A1(KEYINPUT33), .A2(n712), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U785 ( .A(n715), .B(KEYINPUT99), .ZN(n720) );
  XOR2_X1 U786 ( .A(G1981), .B(KEYINPUT100), .Z(n716) );
  XNOR2_X1 U787 ( .A(G305), .B(n716), .ZN(n947) );
  NAND2_X1 U788 ( .A1(n958), .A2(KEYINPUT33), .ZN(n717) );
  OR2_X1 U789 ( .A1(n691), .A2(n717), .ZN(n718) );
  AND2_X1 U790 ( .A1(n947), .A2(n718), .ZN(n719) );
  NAND2_X1 U791 ( .A1(G8), .A2(G166), .ZN(n721) );
  NOR2_X1 U792 ( .A1(G2090), .A2(n721), .ZN(n722) );
  XNOR2_X1 U793 ( .A(n722), .B(KEYINPUT101), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U795 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U796 ( .A(n727), .B(KEYINPUT24), .Z(n728) );
  NAND2_X1 U797 ( .A1(G131), .A2(n901), .ZN(n730) );
  NAND2_X1 U798 ( .A1(G107), .A2(n897), .ZN(n729) );
  NAND2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U800 ( .A1(G119), .A2(n898), .ZN(n731) );
  XNOR2_X1 U801 ( .A(KEYINPUT89), .B(n731), .ZN(n732) );
  NOR2_X1 U802 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U803 ( .A1(G95), .A2(n902), .ZN(n734) );
  NAND2_X1 U804 ( .A1(n735), .A2(n734), .ZN(n911) );
  NAND2_X1 U805 ( .A1(G1991), .A2(n911), .ZN(n736) );
  XNOR2_X1 U806 ( .A(n736), .B(KEYINPUT90), .ZN(n745) );
  NAND2_X1 U807 ( .A1(G117), .A2(n897), .ZN(n738) );
  NAND2_X1 U808 ( .A1(G129), .A2(n898), .ZN(n737) );
  NAND2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U810 ( .A1(n902), .A2(G105), .ZN(n739) );
  XOR2_X1 U811 ( .A(KEYINPUT38), .B(n739), .Z(n740) );
  NOR2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U813 ( .A1(n901), .A2(G141), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n914) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n914), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n769) );
  INV_X1 U817 ( .A(n769), .ZN(n979) );
  XOR2_X1 U818 ( .A(G1986), .B(G290), .Z(n945) );
  NAND2_X1 U819 ( .A1(n979), .A2(n945), .ZN(n749) );
  NOR2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n776) );
  NAND2_X1 U821 ( .A1(n749), .A2(n776), .ZN(n761) );
  XNOR2_X1 U822 ( .A(KEYINPUT88), .B(KEYINPUT36), .ZN(n760) );
  NAND2_X1 U823 ( .A1(G140), .A2(n901), .ZN(n751) );
  NAND2_X1 U824 ( .A1(G104), .A2(n902), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U826 ( .A(KEYINPUT34), .B(n752), .ZN(n757) );
  NAND2_X1 U827 ( .A1(G116), .A2(n897), .ZN(n754) );
  NAND2_X1 U828 ( .A1(G128), .A2(n898), .ZN(n753) );
  NAND2_X1 U829 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U830 ( .A(n755), .B(KEYINPUT35), .Z(n756) );
  NOR2_X1 U831 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U832 ( .A(KEYINPUT87), .B(n758), .Z(n759) );
  XNOR2_X1 U833 ( .A(n760), .B(n759), .ZN(n917) );
  XNOR2_X1 U834 ( .A(G2067), .B(KEYINPUT37), .ZN(n774) );
  NOR2_X1 U835 ( .A1(n917), .A2(n774), .ZN(n970) );
  NAND2_X1 U836 ( .A1(n776), .A2(n970), .ZN(n772) );
  NAND2_X1 U837 ( .A1(n761), .A2(n772), .ZN(n762) );
  XNOR2_X1 U838 ( .A(n765), .B(n764), .ZN(n779) );
  NOR2_X1 U839 ( .A1(G1996), .A2(n914), .ZN(n974) );
  NOR2_X1 U840 ( .A1(G1986), .A2(G290), .ZN(n767) );
  NOR2_X1 U841 ( .A1(G1991), .A2(n911), .ZN(n766) );
  XOR2_X1 U842 ( .A(KEYINPUT105), .B(n766), .Z(n977) );
  NOR2_X1 U843 ( .A1(n767), .A2(n977), .ZN(n768) );
  NOR2_X1 U844 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U845 ( .A1(n974), .A2(n770), .ZN(n771) );
  XNOR2_X1 U846 ( .A(n771), .B(KEYINPUT39), .ZN(n773) );
  NAND2_X1 U847 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U848 ( .A1(n917), .A2(n774), .ZN(n972) );
  NAND2_X1 U849 ( .A1(n775), .A2(n972), .ZN(n777) );
  NAND2_X1 U850 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U851 ( .A1(n779), .A2(n778), .ZN(n781) );
  XNOR2_X1 U852 ( .A(n781), .B(n780), .ZN(G329) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  INV_X1 U855 ( .A(G132), .ZN(G219) );
  INV_X1 U856 ( .A(G82), .ZN(G220) );
  NOR2_X1 U857 ( .A1(n783), .A2(n782), .ZN(G160) );
  XOR2_X1 U858 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n785) );
  NAND2_X1 U859 ( .A1(G7), .A2(G661), .ZN(n784) );
  XNOR2_X1 U860 ( .A(n785), .B(n784), .ZN(G223) );
  INV_X1 U861 ( .A(G223), .ZN(n852) );
  NAND2_X1 U862 ( .A1(n852), .A2(G567), .ZN(n786) );
  XOR2_X1 U863 ( .A(KEYINPUT11), .B(n786), .Z(G234) );
  XNOR2_X1 U864 ( .A(G860), .B(KEYINPUT71), .ZN(n791) );
  OR2_X1 U865 ( .A1(n941), .A2(n791), .ZN(G153) );
  NAND2_X1 U866 ( .A1(G868), .A2(G301), .ZN(n788) );
  OR2_X1 U867 ( .A1(n944), .A2(G868), .ZN(n787) );
  NAND2_X1 U868 ( .A1(n788), .A2(n787), .ZN(G284) );
  INV_X1 U869 ( .A(G868), .ZN(n833) );
  NOR2_X1 U870 ( .A1(G286), .A2(n833), .ZN(n790) );
  NOR2_X1 U871 ( .A1(G868), .A2(G299), .ZN(n789) );
  NOR2_X1 U872 ( .A1(n790), .A2(n789), .ZN(G297) );
  NAND2_X1 U873 ( .A1(n791), .A2(G559), .ZN(n792) );
  NAND2_X1 U874 ( .A1(n792), .A2(n944), .ZN(n793) );
  XNOR2_X1 U875 ( .A(n793), .B(KEYINPUT16), .ZN(n794) );
  XNOR2_X1 U876 ( .A(KEYINPUT74), .B(n794), .ZN(G148) );
  NOR2_X1 U877 ( .A1(G868), .A2(n941), .ZN(n795) );
  XOR2_X1 U878 ( .A(KEYINPUT75), .B(n795), .Z(n798) );
  NAND2_X1 U879 ( .A1(G868), .A2(n944), .ZN(n796) );
  NOR2_X1 U880 ( .A1(G559), .A2(n796), .ZN(n797) );
  NOR2_X1 U881 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U882 ( .A(KEYINPUT76), .B(n799), .ZN(G282) );
  NAND2_X1 U883 ( .A1(G111), .A2(n897), .ZN(n806) );
  NAND2_X1 U884 ( .A1(G135), .A2(n901), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G99), .A2(n902), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U887 ( .A1(n898), .A2(G123), .ZN(n802) );
  XOR2_X1 U888 ( .A(KEYINPUT18), .B(n802), .Z(n803) );
  NOR2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n807), .B(KEYINPUT77), .ZN(n976) );
  XNOR2_X1 U892 ( .A(G2096), .B(n976), .ZN(n809) );
  INV_X1 U893 ( .A(G2100), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n809), .A2(n808), .ZN(G156) );
  NAND2_X1 U895 ( .A1(G80), .A2(n810), .ZN(n813) );
  NAND2_X1 U896 ( .A1(G67), .A2(n811), .ZN(n812) );
  NAND2_X1 U897 ( .A1(n813), .A2(n812), .ZN(n817) );
  NAND2_X1 U898 ( .A1(n814), .A2(G93), .ZN(n815) );
  XOR2_X1 U899 ( .A(KEYINPUT78), .B(n815), .Z(n816) );
  NOR2_X1 U900 ( .A1(n817), .A2(n816), .ZN(n820) );
  NAND2_X1 U901 ( .A1(n818), .A2(G55), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n820), .A2(n819), .ZN(n834) );
  NAND2_X1 U903 ( .A1(n944), .A2(G559), .ZN(n831) );
  XNOR2_X1 U904 ( .A(n941), .B(n831), .ZN(n821) );
  NOR2_X1 U905 ( .A1(G860), .A2(n821), .ZN(n822) );
  XOR2_X1 U906 ( .A(n834), .B(n822), .Z(G145) );
  XOR2_X1 U907 ( .A(n941), .B(G299), .Z(n826) );
  XOR2_X1 U908 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n824) );
  XNOR2_X1 U909 ( .A(G166), .B(KEYINPUT83), .ZN(n823) );
  XNOR2_X1 U910 ( .A(n824), .B(n823), .ZN(n825) );
  XNOR2_X1 U911 ( .A(n826), .B(n825), .ZN(n828) );
  XNOR2_X1 U912 ( .A(G290), .B(G288), .ZN(n827) );
  XNOR2_X1 U913 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U914 ( .A(n829), .B(G305), .ZN(n830) );
  XNOR2_X1 U915 ( .A(n830), .B(n834), .ZN(n921) );
  XOR2_X1 U916 ( .A(n921), .B(n831), .Z(n832) );
  NAND2_X1 U917 ( .A1(G868), .A2(n832), .ZN(n836) );
  NAND2_X1 U918 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U919 ( .A1(n836), .A2(n835), .ZN(G295) );
  NAND2_X1 U920 ( .A1(G2084), .A2(G2078), .ZN(n839) );
  XNOR2_X1 U921 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n837) );
  XNOR2_X1 U922 ( .A(n837), .B(KEYINPUT85), .ZN(n838) );
  XNOR2_X1 U923 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U924 ( .A1(n840), .A2(G2090), .ZN(n841) );
  XNOR2_X1 U925 ( .A(KEYINPUT21), .B(n841), .ZN(n842) );
  NAND2_X1 U926 ( .A1(n842), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U927 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U928 ( .A1(G220), .A2(G219), .ZN(n843) );
  XOR2_X1 U929 ( .A(KEYINPUT22), .B(n843), .Z(n844) );
  NOR2_X1 U930 ( .A1(G218), .A2(n844), .ZN(n845) );
  NAND2_X1 U931 ( .A1(G96), .A2(n845), .ZN(n856) );
  NAND2_X1 U932 ( .A1(n856), .A2(G2106), .ZN(n849) );
  NAND2_X1 U933 ( .A1(G69), .A2(G120), .ZN(n846) );
  NOR2_X1 U934 ( .A1(G237), .A2(n846), .ZN(n847) );
  NAND2_X1 U935 ( .A1(G108), .A2(n847), .ZN(n857) );
  NAND2_X1 U936 ( .A1(n857), .A2(G567), .ZN(n848) );
  NAND2_X1 U937 ( .A1(n849), .A2(n848), .ZN(n858) );
  NAND2_X1 U938 ( .A1(G661), .A2(G483), .ZN(n850) );
  XNOR2_X1 U939 ( .A(KEYINPUT86), .B(n850), .ZN(n851) );
  NOR2_X1 U940 ( .A1(n858), .A2(n851), .ZN(n855) );
  NAND2_X1 U941 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n852), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n853) );
  NAND2_X1 U944 ( .A1(G661), .A2(n853), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U946 ( .A1(n855), .A2(n854), .ZN(G188) );
  XOR2_X1 U947 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G69), .ZN(G235) );
  NOR2_X1 U951 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  INV_X1 U953 ( .A(n858), .ZN(G319) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2090), .Z(n860) );
  XNOR2_X1 U955 ( .A(G2072), .B(G2084), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U957 ( .A(n861), .B(G2096), .Z(n863) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2078), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2678), .Z(n865) );
  XNOR2_X1 U961 ( .A(KEYINPUT109), .B(G2100), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(n867), .B(n866), .Z(G227) );
  XNOR2_X1 U964 ( .A(G1991), .B(G2474), .ZN(n877) );
  XOR2_X1 U965 ( .A(G1961), .B(G1981), .Z(n869) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1986), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U968 ( .A(G1971), .B(G1956), .Z(n871) );
  XNOR2_X1 U969 ( .A(G1976), .B(G1966), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U971 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U972 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(G229) );
  NAND2_X1 U975 ( .A1(G100), .A2(n902), .ZN(n878) );
  XOR2_X1 U976 ( .A(KEYINPUT111), .B(n878), .Z(n880) );
  NAND2_X1 U977 ( .A1(n897), .A2(G112), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(KEYINPUT112), .B(n881), .ZN(n886) );
  NAND2_X1 U980 ( .A1(G124), .A2(n898), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(KEYINPUT44), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n901), .A2(G136), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(G162) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n896) );
  NAND2_X1 U986 ( .A1(G139), .A2(n901), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G103), .A2(n902), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n898), .A2(G127), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n889), .B(KEYINPUT114), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G115), .A2(n897), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n966) );
  XNOR2_X1 U995 ( .A(G164), .B(n966), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n913) );
  NAND2_X1 U997 ( .A1(G118), .A2(n897), .ZN(n900) );
  NAND2_X1 U998 ( .A1(G130), .A2(n898), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n901), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n902), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT45), .B(n905), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT113), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n976), .B(n909), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(n914), .B(G162), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n916), .B(n915), .ZN(n919) );
  XNOR2_X1 U1011 ( .A(n917), .B(G160), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n920), .ZN(G395) );
  XNOR2_X1 U1014 ( .A(n944), .B(G286), .ZN(n922) );
  XNOR2_X1 U1015 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1016 ( .A(n923), .B(G171), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n924), .ZN(G397) );
  XOR2_X1 U1018 ( .A(G2454), .B(G2435), .Z(n926) );
  XNOR2_X1 U1019 ( .A(G2438), .B(G2427), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n926), .B(n925), .ZN(n933) );
  XOR2_X1 U1021 ( .A(KEYINPUT107), .B(G2446), .Z(n928) );
  XNOR2_X1 U1022 ( .A(G2443), .B(G2430), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1024 ( .A(n929), .B(G2451), .Z(n931) );
  XNOR2_X1 U1025 ( .A(G1341), .B(G1348), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n931), .B(n930), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(n933), .B(n932), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n934), .A2(G14), .ZN(n940) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n940), .ZN(n937) );
  NOR2_X1 U1030 ( .A1(G227), .A2(G229), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(KEYINPUT49), .B(n935), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(G225) );
  INV_X1 U1035 ( .A(G225), .ZN(G308) );
  INV_X1 U1036 ( .A(G108), .ZN(G238) );
  INV_X1 U1037 ( .A(n940), .ZN(G401) );
  XNOR2_X1 U1038 ( .A(G301), .B(G1961), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n941), .B(G1341), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(n944), .B(G1348), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G168), .B(G1966), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n949), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n963) );
  XNOR2_X1 U1048 ( .A(G166), .B(G1971), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G1956), .B(KEYINPUT121), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n954), .B(G299), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT122), .B(n961), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .Z(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n1046) );
  XNOR2_X1 U1058 ( .A(KEYINPUT55), .B(KEYINPUT116), .ZN(n1037) );
  XOR2_X1 U1059 ( .A(G2072), .B(n966), .Z(n968) );
  XOR2_X1 U1060 ( .A(G164), .B(G2078), .Z(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT50), .B(n969), .Z(n988) );
  INV_X1 U1063 ( .A(n970), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n985) );
  XOR2_X1 U1065 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT51), .B(n975), .Z(n983) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n981) );
  XOR2_X1 U1070 ( .A(G160), .B(G2084), .Z(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(KEYINPUT115), .B(n986), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1076 ( .A(KEYINPUT52), .B(n989), .Z(n990) );
  NOR2_X1 U1077 ( .A1(n1037), .A2(n990), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(KEYINPUT117), .B(n991), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n992), .A2(G29), .ZN(n1044) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n993), .B(G4), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G1956), .B(G20), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G19), .B(G1341), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1086 ( .A(KEYINPUT123), .B(G1981), .Z(n998) );
  XNOR2_X1 U1087 ( .A(G6), .B(n998), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(n1001), .B(KEYINPUT124), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G21), .B(G1966), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1005), .Z(n1013) );
  XNOR2_X1 U1094 ( .A(G1976), .B(G23), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G1971), .B(G22), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1098 ( .A(G1986), .B(G24), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G5), .B(G1961), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1016), .Z(n1017) );
  NOR2_X1 U1105 ( .A1(G16), .A2(n1017), .ZN(n1042) );
  XOR2_X1 U1106 ( .A(G29), .B(KEYINPUT120), .Z(n1039) );
  XNOR2_X1 U1107 ( .A(G1996), .B(G32), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(G1991), .B(G25), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(G2067), .B(G26), .Z(n1020) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(G28), .ZN(n1023) );
  XNOR2_X1 U1112 ( .A(KEYINPUT118), .B(G2072), .ZN(n1021) );
  XNOR2_X1 U1113 ( .A(G33), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1115 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(G27), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1118 ( .A(KEYINPUT53), .B(n1029), .Z(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n1030) );
  XNOR2_X1 U1120 ( .A(n1030), .B(G34), .ZN(n1031) );
  XNOR2_X1 U1121 ( .A(G2084), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1035) );
  XNOR2_X1 U1123 ( .A(G35), .B(G2090), .ZN(n1034) );
  NOR2_X1 U1124 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1125 ( .A(n1037), .B(n1036), .ZN(n1038) );
  NAND2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1127 ( .A1(G11), .A2(n1040), .ZN(n1041) );
  NOR2_X1 U1128 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1129 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NOR2_X1 U1130 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XOR2_X1 U1131 ( .A(KEYINPUT62), .B(n1047), .Z(n1048) );
  XNOR2_X1 U1132 ( .A(KEYINPUT127), .B(n1048), .ZN(G311) );
  INV_X1 U1133 ( .A(G311), .ZN(G150) );
endmodule

