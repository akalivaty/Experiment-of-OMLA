

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  XNOR2_X1 U323 ( .A(n520), .B(KEYINPUT122), .ZN(n291) );
  XNOR2_X1 U324 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U325 ( .A(n353), .B(n313), .ZN(n316) );
  INV_X1 U326 ( .A(KEYINPUT11), .ZN(n323) );
  XNOR2_X1 U327 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U328 ( .A(n326), .B(n325), .ZN(n330) );
  XNOR2_X1 U329 ( .A(n455), .B(KEYINPUT125), .ZN(n589) );
  XOR2_X1 U330 ( .A(KEYINPUT28), .B(n560), .Z(n532) );
  XNOR2_X1 U331 ( .A(n457), .B(G218GAT), .ZN(n458) );
  XNOR2_X1 U332 ( .A(n459), .B(n458), .ZN(G1355GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT97), .B(KEYINPUT4), .Z(n293) );
  XNOR2_X1 U334 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n303) );
  XOR2_X1 U336 ( .A(G1GAT), .B(G127GAT), .Z(n337) );
  XOR2_X1 U337 ( .A(G85GAT), .B(n337), .Z(n295) );
  XOR2_X1 U338 ( .A(G120GAT), .B(G57GAT), .Z(n376) );
  XNOR2_X1 U339 ( .A(G162GAT), .B(n376), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U341 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n297) );
  NAND2_X1 U342 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n299), .B(n298), .Z(n301) );
  XOR2_X1 U345 ( .A(G113GAT), .B(KEYINPUT0), .Z(n414) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G134GAT), .Z(n312) );
  XNOR2_X1 U347 ( .A(n414), .B(n312), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT94), .B(G148GAT), .Z(n305) );
  XNOR2_X1 U351 ( .A(G141GAT), .B(G155GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n307) );
  XOR2_X1 U353 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n306) );
  XOR2_X1 U354 ( .A(n307), .B(n306), .Z(n441) );
  XOR2_X1 U355 ( .A(n308), .B(n441), .Z(n477) );
  XNOR2_X1 U356 ( .A(KEYINPUT99), .B(n477), .ZN(n518) );
  XOR2_X1 U357 ( .A(G43GAT), .B(KEYINPUT7), .Z(n310) );
  XNOR2_X1 U358 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n353) );
  AND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n311) );
  INV_X1 U361 ( .A(n316), .ZN(n315) );
  INV_X1 U362 ( .A(KEYINPUT65), .ZN(n314) );
  NAND2_X1 U363 ( .A1(n315), .A2(n314), .ZN(n318) );
  NAND2_X1 U364 ( .A1(n316), .A2(KEYINPUT65), .ZN(n317) );
  NAND2_X1 U365 ( .A1(n318), .A2(n317), .ZN(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT73), .B(G85GAT), .Z(n320) );
  XNOR2_X1 U367 ( .A(G99GAT), .B(G106GAT), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n372) );
  XOR2_X1 U369 ( .A(n372), .B(KEYINPUT10), .Z(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U371 ( .A(G50GAT), .B(G162GAT), .Z(n446) );
  XNOR2_X1 U372 ( .A(n446), .B(KEYINPUT9), .ZN(n324) );
  XOR2_X1 U373 ( .A(G92GAT), .B(KEYINPUT77), .Z(n328) );
  XNOR2_X1 U374 ( .A(G190GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U375 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U376 ( .A(G36GAT), .B(n329), .Z(n400) );
  XOR2_X1 U377 ( .A(n330), .B(n400), .Z(n557) );
  XNOR2_X1 U378 ( .A(n557), .B(KEYINPUT78), .ZN(n577) );
  XNOR2_X1 U379 ( .A(KEYINPUT36), .B(n577), .ZN(n493) );
  XOR2_X1 U380 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n332) );
  XNOR2_X1 U381 ( .A(G57GAT), .B(G64GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U383 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n334) );
  XNOR2_X1 U384 ( .A(KEYINPUT15), .B(KEYINPUT82), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n349) );
  XOR2_X1 U387 ( .A(G71GAT), .B(KEYINPUT13), .Z(n375) );
  XOR2_X1 U388 ( .A(n375), .B(n337), .Z(n339) );
  XNOR2_X1 U389 ( .A(G211GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n345) );
  XOR2_X1 U391 ( .A(G8GAT), .B(KEYINPUT69), .Z(n341) );
  XNOR2_X1 U392 ( .A(G15GAT), .B(G22GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n352) );
  XOR2_X1 U394 ( .A(KEYINPUT14), .B(n352), .Z(n343) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(n345), .B(n344), .Z(n347) );
  XNOR2_X1 U398 ( .A(G183GAT), .B(G155GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n588) );
  INV_X1 U401 ( .A(n588), .ZN(n574) );
  NOR2_X1 U402 ( .A1(n493), .A2(n574), .ZN(n351) );
  XNOR2_X1 U403 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n387) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n366) );
  XOR2_X1 U406 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n355) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U409 ( .A(n356), .B(KEYINPUT67), .Z(n364) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G36GAT), .Z(n358) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(G50GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U413 ( .A(G1GAT), .B(G197GAT), .Z(n360) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G141GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n564) );
  INV_X1 U419 ( .A(n564), .ZN(n583) );
  XOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n368) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U423 ( .A(n369), .B(KEYINPUT70), .Z(n374) );
  XOR2_X1 U424 ( .A(KEYINPUT75), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G204GAT), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n397) );
  XNOR2_X1 U427 ( .A(n372), .B(n397), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n380) );
  XOR2_X1 U429 ( .A(n375), .B(G92GAT), .Z(n378) );
  XNOR2_X1 U430 ( .A(G148GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n385) );
  XOR2_X1 U433 ( .A(KEYINPUT72), .B(G78GAT), .Z(n436) );
  XOR2_X1 U434 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n382) );
  XNOR2_X1 U435 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n436), .B(n383), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n465) );
  INV_X1 U439 ( .A(n465), .ZN(n460) );
  NOR2_X1 U440 ( .A1(n583), .A2(n460), .ZN(n386) );
  NAND2_X1 U441 ( .A1(n387), .A2(n386), .ZN(n395) );
  XOR2_X1 U442 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n393) );
  XNOR2_X1 U443 ( .A(n465), .B(KEYINPUT64), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n388), .B(KEYINPUT41), .ZN(n567) );
  NAND2_X1 U445 ( .A1(n567), .A2(n583), .ZN(n389) );
  XOR2_X1 U446 ( .A(KEYINPUT46), .B(n389), .Z(n390) );
  NOR2_X1 U447 ( .A1(n588), .A2(n390), .ZN(n391) );
  NAND2_X1 U448 ( .A1(n391), .A2(n557), .ZN(n392) );
  XOR2_X1 U449 ( .A(n393), .B(n392), .Z(n394) );
  AND2_X1 U450 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT48), .B(n396), .ZN(n528) );
  INV_X1 U452 ( .A(n528), .ZN(n411) );
  XOR2_X1 U453 ( .A(n397), .B(KEYINPUT100), .Z(n399) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U456 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U457 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT92), .B(G211GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(n404), .ZN(n451) );
  XOR2_X1 U461 ( .A(G8GAT), .B(n451), .Z(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U463 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U466 ( .A(G169GAT), .B(n409), .Z(n430) );
  XNOR2_X1 U467 ( .A(n410), .B(n430), .ZN(n520) );
  NAND2_X1 U468 ( .A1(n411), .A2(n291), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n412), .B(KEYINPUT54), .ZN(n413) );
  NOR2_X1 U470 ( .A1(n518), .A2(n413), .ZN(n561) );
  XOR2_X1 U471 ( .A(n414), .B(G120GAT), .Z(n416) );
  NAND2_X1 U472 ( .A1(G227GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U474 ( .A(n417), .B(G99GAT), .Z(n422) );
  XOR2_X1 U475 ( .A(G176GAT), .B(KEYINPUT20), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U478 ( .A(G43GAT), .B(n420), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U480 ( .A(G71GAT), .B(G190GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(G15GAT), .B(G134GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n432) );
  XOR2_X1 U484 ( .A(KEYINPUT88), .B(KEYINPUT84), .Z(n428) );
  XNOR2_X1 U485 ( .A(G127GAT), .B(KEYINPUT85), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n563) );
  XOR2_X1 U489 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n434) );
  XNOR2_X1 U490 ( .A(G218GAT), .B(G106GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U492 ( .A(n435), .B(KEYINPUT96), .Z(n438) );
  XNOR2_X1 U493 ( .A(G22GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n450) );
  XOR2_X1 U495 ( .A(KEYINPUT89), .B(KEYINPUT95), .Z(n440) );
  XNOR2_X1 U496 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U498 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n444) );
  NAND2_X1 U500 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n560) );
  NOR2_X1 U506 ( .A1(n563), .A2(n560), .ZN(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT26), .B(KEYINPUT102), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n547) );
  NAND2_X1 U509 ( .A1(n561), .A2(n547), .ZN(n455) );
  INV_X1 U510 ( .A(n589), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n456), .A2(n493), .ZN(n459) );
  INV_X1 U512 ( .A(KEYINPUT62), .ZN(n457) );
  INV_X1 U513 ( .A(G204GAT), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n462) );
  NAND2_X1 U515 ( .A1(n589), .A2(n460), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(G1353GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n483) );
  NAND2_X1 U519 ( .A1(n465), .A2(n583), .ZN(n495) );
  NAND2_X1 U520 ( .A1(n577), .A2(n588), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT83), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT16), .B(n467), .ZN(n481) );
  INV_X1 U523 ( .A(n563), .ZN(n576) );
  XNOR2_X1 U524 ( .A(n520), .B(KEYINPUT27), .ZN(n473) );
  NAND2_X1 U525 ( .A1(n518), .A2(n473), .ZN(n529) );
  NOR2_X1 U526 ( .A1(n529), .A2(n532), .ZN(n468) );
  XOR2_X1 U527 ( .A(KEYINPUT101), .B(n468), .Z(n469) );
  NAND2_X1 U528 ( .A1(n576), .A2(n469), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n520), .A2(n563), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n470), .A2(n560), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT25), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT103), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n473), .A2(n547), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n480), .B(KEYINPUT104), .ZN(n491) );
  NAND2_X1 U538 ( .A1(n481), .A2(n491), .ZN(n505) );
  NOR2_X1 U539 ( .A1(n495), .A2(n505), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n488), .A2(n518), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n520), .A2(n488), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U546 ( .A1(n488), .A2(n563), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n532), .A2(n488), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT106), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n574), .ZN(n492) );
  NOR2_X1 U552 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n494), .ZN(n515) );
  NOR2_X1 U554 ( .A1(n515), .A2(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(n496), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n518), .A2(n503), .ZN(n498) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n503), .A2(n520), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n501) );
  NAND2_X1 U562 ( .A1(n563), .A2(n503), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n532), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  NAND2_X1 U568 ( .A1(n564), .A2(n567), .ZN(n516) );
  NOR2_X1 U569 ( .A1(n516), .A2(n505), .ZN(n511) );
  NAND2_X1 U570 ( .A1(n518), .A2(n511), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n520), .A2(n511), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n563), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n532), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT110), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n518), .A2(n524), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n524), .A2(n520), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U588 ( .A1(n563), .A2(n524), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n526) );
  NAND2_X1 U591 ( .A1(n524), .A2(n532), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n534) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT114), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n563), .A2(n548), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n544), .A2(n583), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U603 ( .A1(n544), .A2(n567), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U605 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n540) );
  NAND2_X1 U608 ( .A1(n544), .A2(n588), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  INV_X1 U612 ( .A(n577), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT120), .B(n549), .Z(n555) );
  NAND2_X1 U617 ( .A1(n555), .A2(n583), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U620 ( .A1(n567), .A2(n555), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n555), .A2(n588), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n559) );
  INV_X1 U626 ( .A(n555), .ZN(n556) );
  NOR2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(KEYINPUT55), .B(n562), .ZN(n579) );
  NAND2_X1 U631 ( .A1(n579), .A2(n563), .ZN(n573) );
  NOR2_X1 U632 ( .A1(n564), .A2(n573), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  INV_X1 U635 ( .A(n567), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n568), .A2(n576), .ZN(n569) );
  AND2_X1 U637 ( .A1(n579), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(n572), .ZN(G1349GAT) );
  NOR2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(G183GAT), .B(n575), .Z(G1350GAT) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  AND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n582), .B(G190GAT), .Z(G1351GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n589), .ZN(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n585) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1352GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
endmodule

