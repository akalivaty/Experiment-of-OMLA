//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(new_n189), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(KEYINPUT1), .B2(new_n189), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n191), .A2(new_n194), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT84), .B1(new_n198), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT10), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT84), .B(KEYINPUT10), .C1(new_n198), .C2(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n217), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n206), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n223), .A3(G101), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n195), .A2(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n192), .A2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n229), .B1(new_n232), .B2(new_n188), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n229), .B(new_n235), .C1(new_n232), .C2(new_n188), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n225), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n222), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .A3(KEYINPUT11), .A4(G134), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT11), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(G137), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n243), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G131), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(G131), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n244), .A2(new_n245), .B1(new_n240), .B2(G137), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n241), .A4(new_n243), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n215), .A2(new_n238), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n191), .A2(new_n194), .A3(new_n197), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(new_n210), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n198), .A2(new_n210), .ZN(new_n261));
  INV_X1    g075(.A(new_n210), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT12), .B(new_n253), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n255), .A2(new_n256), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n256), .B1(new_n255), .B2(new_n265), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XNOR2_X1  g087(.A(G110), .B(G140), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n266), .A2(new_n267), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n215), .A2(new_n238), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n253), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n255), .A3(new_n275), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT86), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n267), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n255), .A2(new_n256), .A3(new_n265), .ZN(new_n283));
  INV_X1    g097(.A(new_n275), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT86), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n279), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n187), .B(G469), .C1(new_n288), .C2(G902), .ZN(new_n289));
  INV_X1    g103(.A(G221), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT9), .B(G234), .Z(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G475), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT18), .A2(G131), .ZN(new_n297));
  INV_X1    g111(.A(G237), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n272), .A2(G214), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n192), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n272), .A2(G143), .A3(G214), .A4(new_n298), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n297), .B1(new_n302), .B2(KEYINPUT92), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(KEYINPUT92), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(new_n195), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(KEYINPUT92), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  OR3_X1    g125(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n195), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(G146), .A3(new_n312), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n250), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n302), .A2(KEYINPUT17), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n302), .A2(new_n317), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n300), .A2(new_n250), .A3(new_n301), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n316), .B(new_n318), .C1(new_n321), .C2(KEYINPUT17), .ZN(new_n322));
  XNOR2_X1  g136(.A(G113), .B(G122), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(new_n199), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT94), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n309), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n306), .B(KEYINPUT19), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n195), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n328), .A2(KEYINPUT93), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(KEYINPUT93), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n321), .A2(new_n329), .A3(new_n315), .A4(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n324), .B1(new_n309), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n296), .B(new_n292), .C1(new_n326), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT95), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n309), .A2(new_n322), .A3(new_n325), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n309), .A2(new_n331), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n324), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT95), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n296), .A4(new_n292), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT20), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n324), .B1(new_n309), .B2(new_n322), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n292), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G475), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n333), .A2(KEYINPUT95), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n268), .A2(G952), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(G234), .B2(G237), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT21), .B(G898), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n349), .B(KEYINPUT97), .Z(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(new_n292), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G128), .B(G143), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(new_n240), .ZN(new_n355));
  INV_X1    g169(.A(G116), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT14), .A3(G122), .ZN(new_n357));
  XNOR2_X1  g171(.A(G116), .B(G122), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(G107), .B(new_n357), .C1(new_n359), .C2(KEYINPUT14), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n355), .B(new_n360), .C1(G107), .C2(new_n359), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n192), .A2(G128), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n362), .B(G134), .C1(KEYINPUT13), .C2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n358), .B(new_n202), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n354), .A2(new_n240), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n291), .A2(G217), .A3(new_n268), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n292), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT15), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n372), .A2(KEYINPUT96), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(KEYINPUT96), .ZN(new_n374));
  OAI21_X1  g188(.A(G478), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n371), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n346), .A2(new_n353), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G214), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G119), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n356), .A2(G119), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT2), .B(G113), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G113), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT2), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G113), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n384), .A2(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n224), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT89), .B1(new_n222), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n396), .B(new_n393), .C1(new_n220), .C2(new_n221), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(G110), .B(G122), .Z(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT5), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(G113), .C1(KEYINPUT5), .C2(new_n382), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n384), .B2(new_n385), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n210), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n233), .A2(G125), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n198), .B2(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n268), .A2(G224), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT7), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n408), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n403), .B(new_n262), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n399), .B(KEYINPUT8), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n406), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n292), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n222), .A2(new_n394), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n396), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n222), .A2(new_n394), .A3(KEYINPUT89), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n405), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n399), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT90), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n419), .A2(new_n423), .A3(new_n420), .A4(new_n399), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n399), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n395), .A2(new_n397), .A3(new_n404), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n420), .B1(new_n426), .B2(new_n400), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n422), .A2(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n409), .B(KEYINPUT91), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n408), .B(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n415), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G210), .B1(G237), .B2(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(new_n406), .A3(KEYINPUT6), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n400), .B1(new_n398), .B2(new_n405), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n423), .B1(new_n435), .B2(new_n420), .ZN(new_n436));
  INV_X1    g250(.A(new_n424), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n430), .B(new_n434), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n414), .A2(new_n292), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n432), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n380), .B1(new_n433), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G469), .B1(new_n288), .B2(G902), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n278), .A2(new_n255), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n284), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(KEYINPUT88), .A3(new_n284), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n255), .A2(new_n265), .A3(new_n275), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n292), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n444), .A2(KEYINPUT87), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n295), .A2(new_n378), .A3(new_n443), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n234), .A2(new_n236), .B1(new_n252), .B2(new_n249), .ZN(new_n457));
  OR3_X1    g271(.A1(new_n240), .A2(KEYINPUT66), .A3(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n240), .A2(G137), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n458), .B(G131), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n258), .A2(new_n252), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n456), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n236), .ZN(new_n464));
  OAI22_X1  g278(.A1(new_n193), .A2(new_n196), .B1(new_n230), .B2(new_n231), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n235), .B1(new_n465), .B2(new_n229), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n253), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n258), .A2(new_n252), .A3(new_n461), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT72), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n387), .A2(new_n392), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(KEYINPUT73), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(new_n470), .A3(new_n468), .ZN(new_n477));
  INV_X1    g291(.A(new_n470), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n249), .A2(new_n252), .B1(new_n465), .B2(new_n229), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n462), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n272), .A2(G210), .A3(new_n298), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(G101), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT71), .ZN(new_n489));
  OR3_X1    g303(.A1(new_n483), .A2(KEYINPUT29), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n471), .A2(KEYINPUT73), .A3(new_n472), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT73), .B1(new_n471), .B2(new_n472), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n488), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n467), .A2(new_n468), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n478), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n477), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT29), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n462), .B2(new_n479), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n502), .B(new_n478), .C1(new_n495), .C2(new_n501), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n477), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n488), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n490), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n292), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G472), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n494), .A2(new_n503), .A3(new_n477), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n494), .A2(new_n503), .A3(KEYINPUT31), .A4(new_n477), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n491), .A2(new_n492), .A3(new_n481), .ZN(new_n515));
  INV_X1    g329(.A(new_n489), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT74), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n483), .A2(new_n489), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT74), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n514), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT75), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n509), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT32), .B(new_n524), .C1(new_n518), .C2(new_n521), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n508), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT79), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n530), .B(new_n531), .Z(new_n532));
  NAND2_X1  g346(.A1(new_n381), .A2(G128), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n189), .A2(G119), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT24), .B(G110), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT77), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n314), .A2(new_n315), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n533), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G110), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(new_n546), .A3(new_n538), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n540), .A2(new_n541), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n306), .A2(new_n195), .ZN(new_n549));
  OAI22_X1  g363(.A1(new_n536), .A2(new_n538), .B1(G110), .B2(new_n544), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n315), .B(new_n549), .C1(new_n550), .C2(KEYINPUT78), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n532), .B1(new_n553), .B2(KEYINPUT80), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(KEYINPUT80), .B2(new_n553), .ZN(new_n555));
  INV_X1    g369(.A(new_n553), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n532), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n559), .A2(new_n292), .B1(KEYINPUT81), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n562));
  AOI211_X1 g376(.A(G902), .B(new_n562), .C1(new_n555), .C2(new_n558), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G217), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(new_n292), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G902), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT82), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n564), .A2(new_n566), .B1(new_n568), .B2(new_n559), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n528), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n455), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n204), .ZN(G3));
  AND3_X1   g386(.A1(new_n519), .A2(new_n520), .A3(new_n514), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n520), .B1(new_n519), .B2(new_n514), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n292), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(G472), .B1(new_n522), .B2(new_n525), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n295), .A2(new_n569), .A3(new_n454), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT99), .B1(new_n578), .B2(new_n380), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n379), .C1(new_n431), .C2(new_n432), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n380), .A2(KEYINPUT98), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n431), .B2(new_n432), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n581), .ZN(new_n586));
  INV_X1    g400(.A(new_n584), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n577), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n370), .B1(KEYINPUT100), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(KEYINPUT100), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(G478), .A3(new_n292), .ZN(new_n594));
  AOI21_X1  g408(.A(G478), .B1(new_n370), .B2(new_n292), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT101), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n346), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n353), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT34), .B(G104), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NOR3_X1   g416(.A1(new_n346), .A2(new_n353), .A3(new_n376), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n589), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NOR2_X1   g420(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n553), .B(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n564), .A2(new_n566), .B1(new_n568), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n576), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n455), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT37), .B(G110), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G12));
  NAND2_X1  g428(.A1(new_n295), .A2(new_n454), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n525), .B1(new_n573), .B2(new_n574), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT32), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n522), .A2(new_n509), .A3(new_n525), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n617), .A2(new_n618), .B1(G472), .B2(new_n507), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n609), .B1(new_n588), .B2(new_n585), .ZN(new_n621));
  INV_X1    g435(.A(new_n346), .ZN(new_n622));
  INV_X1    g436(.A(new_n348), .ZN(new_n623));
  INV_X1    g437(.A(new_n352), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(G900), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n622), .A2(new_n377), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  NAND2_X1  g442(.A1(new_n433), .A2(new_n442), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n346), .A2(new_n377), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n625), .B(KEYINPUT39), .Z(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n295), .A2(new_n454), .A3(new_n634), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n610), .B(new_n632), .C1(new_n635), .C2(KEYINPUT40), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n617), .A2(new_n618), .ZN(new_n637));
  INV_X1    g451(.A(new_n510), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n489), .A2(new_n497), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n639), .B2(KEYINPUT103), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(KEYINPUT103), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n292), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n635), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n380), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n631), .A2(new_n636), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT104), .B(G143), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G45));
  AND3_X1   g464(.A1(new_n597), .A2(new_n346), .A3(new_n625), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n620), .A2(new_n621), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  NAND2_X1  g467(.A1(new_n451), .A2(new_n292), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G469), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n453), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n293), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n584), .B1(new_n579), .B2(new_n581), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n528), .A2(new_n569), .A3(new_n599), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT41), .B(G113), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  NAND3_X1  g478(.A1(new_n528), .A2(new_n569), .A3(new_n603), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n356), .ZN(G18));
  OAI211_X1 g481(.A(new_n610), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n528), .A2(new_n378), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n381), .ZN(G21));
  AOI21_X1  g485(.A(G902), .B1(new_n518), .B2(new_n521), .ZN(new_n672));
  INV_X1    g486(.A(G472), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT106), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n575), .A2(new_n675), .A3(G472), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n524), .B(KEYINPUT105), .Z(new_n677));
  AOI21_X1  g491(.A(new_n516), .B1(new_n493), .B2(new_n498), .ZN(new_n678));
  INV_X1    g492(.A(new_n514), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n674), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n353), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n569), .A3(new_n682), .A4(new_n657), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n377), .B(new_n346), .C1(new_n658), .C2(new_n659), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT107), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n569), .A2(new_n674), .A3(new_n676), .A4(new_n680), .ZN(new_n686));
  INV_X1    g500(.A(new_n657), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(new_n353), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n632), .B1(new_n588), .B2(new_n585), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT108), .B(G122), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G24));
  NAND4_X1  g508(.A1(new_n651), .A2(new_n674), .A3(new_n676), .A4(new_n680), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n668), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  AND3_X1   g511(.A1(new_n433), .A2(new_n442), .A3(new_n379), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n452), .A2(new_n292), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n276), .A2(new_n280), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(G469), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n453), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n698), .A2(new_n699), .A3(new_n294), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n578), .A2(new_n380), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n703), .A3(new_n433), .A4(new_n294), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n526), .B2(new_n527), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n617), .A2(KEYINPUT110), .A3(new_n618), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n508), .A3(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n708), .A2(new_n569), .A3(new_n651), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n570), .B1(new_n704), .B2(new_n707), .ZN(new_n715));
  INV_X1    g529(.A(new_n651), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(G131), .Z(G33));
  NAND2_X1  g534(.A1(new_n715), .A2(new_n626), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  INV_X1    g536(.A(new_n698), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n622), .A2(new_n597), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT43), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n576), .A2(new_n609), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(KEYINPUT43), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n452), .B1(new_n701), .B2(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n288), .B2(KEYINPUT45), .ZN(new_n732));
  INV_X1    g546(.A(new_n700), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n453), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT46), .B1(new_n732), .B2(new_n733), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n294), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n633), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n730), .B(new_n738), .C1(new_n729), .C2(new_n728), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  NOR3_X1   g554(.A1(new_n723), .A2(new_n716), .A3(new_n569), .ZN(new_n741));
  NAND2_X1  g555(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n737), .A2(KEYINPUT111), .ZN(new_n743));
  NOR2_X1   g557(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(new_n294), .C1(new_n735), .C2(new_n736), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n742), .A2(new_n743), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n745), .B1(new_n743), .B2(new_n747), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n619), .B(new_n741), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  AND2_X1   g565(.A1(new_n656), .A2(KEYINPUT49), .ZN(new_n752));
  INV_X1    g566(.A(new_n569), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n631), .A2(new_n752), .A3(new_n753), .A4(new_n380), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n294), .B1(new_n656), .B2(KEYINPUT49), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n644), .A2(new_n755), .A3(new_n724), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT113), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n748), .A2(new_n749), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n294), .B2(new_n656), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n725), .A2(new_n727), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n623), .A3(new_n686), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n698), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n657), .A2(new_n698), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n764), .A2(new_n644), .A3(new_n753), .A4(new_n623), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n622), .A3(new_n596), .A4(new_n594), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n761), .A2(new_n623), .A3(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n610), .A3(new_n681), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n631), .A2(new_n379), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n657), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n763), .A2(KEYINPUT51), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n763), .B2(new_n775), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n776), .A2(new_n777), .A3(new_n347), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n660), .B1(new_n661), .B2(new_n665), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n670), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n622), .A2(new_n376), .A3(new_n625), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n615), .A2(new_n619), .A3(new_n723), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n695), .B1(new_n704), .B2(new_n707), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n610), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n692), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n455), .B1(new_n570), .B2(new_n611), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n340), .A2(new_n345), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n377), .A4(new_n343), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT114), .B1(new_n346), .B2(new_n376), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n598), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n682), .A3(new_n443), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n577), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n714), .A2(new_n794), .A3(new_n718), .A4(new_n721), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n644), .A2(new_n609), .A3(new_n703), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n690), .A3(new_n294), .A4(new_n625), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n620), .B(new_n621), .C1(new_n626), .C2(new_n651), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n696), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n696), .A3(new_n798), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT52), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n785), .A2(new_n795), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n800), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n692), .A2(new_n780), .A3(new_n784), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n714), .A2(new_n794), .A3(new_n718), .A4(new_n721), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n810), .A3(new_n811), .A4(KEYINPUT53), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n803), .A2(new_n804), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n805), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n807), .A2(new_n810), .A3(KEYINPUT116), .A4(KEYINPUT53), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n803), .B2(new_n804), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n808), .B2(new_n809), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n821), .A3(new_n807), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n816), .A2(new_n818), .B1(new_n822), .B2(new_n804), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n778), .B(new_n815), .C1(new_n823), .C2(new_n813), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n762), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT118), .Z(new_n826));
  AND3_X1   g640(.A1(new_n765), .A2(new_n346), .A3(new_n597), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n767), .A2(new_n569), .A3(new_n712), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT48), .Z(new_n829));
  NOR4_X1   g643(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(G952), .A2(G953), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n758), .B1(new_n830), .B2(new_n831), .ZN(G75));
  NAND3_X1  g646(.A1(new_n805), .A2(new_n814), .A3(new_n812), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(G210), .A3(G902), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n428), .B(new_n430), .Z(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT55), .Z(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n272), .A2(G952), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n838), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n834), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT119), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n839), .A2(new_n846), .A3(new_n841), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(G51));
  NAND2_X1  g662(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n815), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n700), .B(KEYINPUT57), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n854), .A3(new_n851), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n451), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n732), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n833), .A2(G902), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n840), .B1(new_n856), .B2(new_n858), .ZN(G54));
  NAND4_X1  g673(.A1(new_n833), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n860));
  INV_X1    g674(.A(new_n337), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n840), .ZN(G60));
  NAND2_X1  g678(.A1(G478), .A2(G902), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT59), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n850), .A2(new_n593), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n815), .B1(new_n823), .B2(new_n813), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n593), .B1(new_n868), .B2(new_n866), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n869), .A3(new_n840), .ZN(G63));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n565), .A2(new_n292), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n559), .B1(new_n833), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n840), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n833), .A2(new_n608), .A3(new_n873), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n833), .A2(KEYINPUT122), .A3(new_n608), .A4(new_n873), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(G66));
  AOI21_X1  g696(.A(new_n268), .B1(new_n350), .B2(G224), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n692), .A2(new_n780), .A3(new_n794), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n272), .ZN(new_n885));
  INV_X1    g699(.A(G898), .ZN(new_n886));
  INV_X1    g700(.A(new_n272), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n428), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n885), .B(new_n888), .ZN(G69));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n719), .B1(new_n626), .B2(new_n715), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n696), .A2(new_n798), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n690), .A2(new_n569), .A3(new_n712), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n738), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n750), .A3(new_n739), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n272), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n272), .A2(G900), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n890), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT125), .B(new_n897), .C1(new_n895), .C2(new_n272), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n502), .B1(new_n495), .B2(new_n501), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n327), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n648), .A2(new_n892), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(KEYINPUT62), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n648), .A2(new_n907), .A3(new_n892), .ZN(new_n908));
  INV_X1    g722(.A(new_n570), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n645), .A3(new_n698), .A4(new_n791), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n739), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI221_X1 g728(.A(new_n750), .B1(new_n906), .B2(new_n908), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n904), .B1(new_n915), .B2(new_n272), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT126), .B1(new_n903), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n899), .ZN(new_n918));
  INV_X1    g732(.A(new_n900), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n904), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n750), .B1(new_n914), .B2(new_n912), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n906), .A2(new_n908), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n272), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n902), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(G227), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n897), .B1(new_n927), .B2(new_n887), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n917), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n917), .B2(new_n926), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(G72));
  OR2_X1    g746(.A1(new_n915), .A2(new_n884), .ZN(new_n933));
  NAND2_X1  g747(.A1(G472), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT63), .Z(new_n935));
  AOI21_X1  g749(.A(new_n488), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n840), .B1(new_n936), .B2(new_n504), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n823), .B1(new_n505), .B2(new_n510), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n935), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n935), .B1(new_n895), .B2(new_n884), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT127), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(new_n477), .A3(new_n503), .A4(new_n488), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n937), .A2(new_n939), .A3(new_n942), .ZN(G57));
endmodule


