

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764;

  XNOR2_X1 U369 ( .A(n645), .B(n647), .ZN(n648) );
  BUF_X1 U370 ( .A(n585), .Z(n348) );
  NOR2_X1 U371 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U372 ( .A1(n403), .A2(n522), .ZN(n393) );
  AND2_X1 U373 ( .A1(n408), .A2(n407), .ZN(n350) );
  INV_X1 U374 ( .A(KEYINPUT67), .ZN(n460) );
  NOR2_X2 U375 ( .A1(n652), .A2(n574), .ZN(n571) );
  AND2_X2 U376 ( .A1(n347), .A2(n346), .ZN(n394) );
  INV_X1 U377 ( .A(n398), .ZN(n346) );
  NAND2_X1 U378 ( .A1(n391), .A2(n402), .ZN(n347) );
  OR2_X2 U379 ( .A1(n612), .A2(n526), .ZN(n360) );
  XNOR2_X1 U380 ( .A(n745), .B(n515), .ZN(n644) );
  XNOR2_X2 U381 ( .A(n507), .B(n508), .ZN(n745) );
  XNOR2_X2 U382 ( .A(n478), .B(n405), .ZN(n404) );
  NOR2_X1 U383 ( .A1(G953), .A2(G237), .ZN(n467) );
  XNOR2_X1 U384 ( .A(G101), .B(G104), .ZN(n488) );
  XNOR2_X1 U385 ( .A(n424), .B(G953), .ZN(n755) );
  NAND2_X2 U386 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X2 U387 ( .A(n531), .B(KEYINPUT22), .ZN(n538) );
  NOR2_X2 U388 ( .A1(n369), .A2(n380), .ZN(n531) );
  NAND2_X1 U389 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X1 U390 ( .A1(n631), .A2(n754), .ZN(n692) );
  XNOR2_X1 U391 ( .A(n475), .B(n474), .ZN(n557) );
  XNOR2_X1 U392 ( .A(n388), .B(n443), .ZN(n735) );
  XOR2_X1 U393 ( .A(KEYINPUT59), .B(n639), .Z(n640) );
  XNOR2_X1 U394 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n480) );
  BUF_X1 U395 ( .A(G107), .Z(n374) );
  INV_X1 U396 ( .A(KEYINPUT64), .ZN(n424) );
  XNOR2_X1 U397 ( .A(G902), .B(KEYINPUT15), .ZN(n580) );
  NAND2_X1 U398 ( .A1(n379), .A2(n414), .ZN(n371) );
  NAND2_X2 U399 ( .A1(n379), .A2(n414), .ZN(n376) );
  XNOR2_X2 U400 ( .A(n751), .B(G146), .ZN(n495) );
  XNOR2_X2 U401 ( .A(n404), .B(n513), .ZN(n751) );
  BUF_X1 U402 ( .A(n636), .Z(n349) );
  XNOR2_X1 U403 ( .A(n632), .B(n418), .ZN(n417) );
  NAND2_X1 U404 ( .A1(n699), .A2(n698), .ZN(n695) );
  AND2_X1 U405 ( .A1(n617), .A2(n385), .ZN(n384) );
  NOR2_X1 U406 ( .A1(n685), .A2(n622), .ZN(n385) );
  NAND2_X1 U407 ( .A1(n518), .A2(n580), .ZN(n406) );
  XNOR2_X1 U408 ( .A(n432), .B(n355), .ZN(n698) );
  XNOR2_X1 U409 ( .A(n356), .B(KEYINPUT98), .ZN(n355) );
  INV_X1 U410 ( .A(KEYINPUT21), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n441), .B(n440), .ZN(n448) );
  XNOR2_X1 U412 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n440) );
  XOR2_X1 U413 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n463) );
  INV_X1 U414 ( .A(n415), .ZN(n412) );
  XNOR2_X1 U415 ( .A(n389), .B(KEYINPUT68), .ZN(n603) );
  NAND2_X1 U416 ( .A1(n565), .A2(n390), .ZN(n389) );
  AND2_X1 U417 ( .A1(n592), .A2(n698), .ZN(n390) );
  OR2_X1 U418 ( .A1(n735), .A2(G902), .ZN(n387) );
  XNOR2_X1 U419 ( .A(G119), .B(G137), .ZN(n435) );
  XNOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT24), .ZN(n438) );
  XOR2_X1 U421 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n439) );
  INV_X1 U422 ( .A(KEYINPUT10), .ZN(n433) );
  XNOR2_X1 U423 ( .A(n366), .B(n637), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n638), .B(KEYINPUT91), .ZN(n738) );
  INV_X1 U425 ( .A(KEYINPUT87), .ZN(n549) );
  NAND2_X1 U426 ( .A1(n519), .A2(n627), .ZN(n407) );
  NAND2_X1 U427 ( .A1(n400), .A2(n522), .ZN(n399) );
  XNOR2_X1 U428 ( .A(G116), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X1 U429 ( .A(n383), .B(n382), .ZN(n626) );
  INV_X1 U430 ( .A(KEYINPUT48), .ZN(n382) );
  XNOR2_X1 U431 ( .A(n477), .B(G134), .ZN(n405) );
  AND2_X1 U432 ( .A1(n628), .A2(KEYINPUT65), .ZN(n415) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n421) );
  INV_X1 U434 ( .A(G237), .ZN(n498) );
  INV_X1 U435 ( .A(G902), .ZN(n499) );
  INV_X1 U436 ( .A(G953), .ZN(n739) );
  XOR2_X1 U437 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n452) );
  XNOR2_X1 U438 ( .A(KEYINPUT104), .B(KEYINPUT106), .ZN(n451) );
  NAND2_X1 U439 ( .A1(n448), .A2(G217), .ZN(n450) );
  XNOR2_X1 U440 ( .A(G134), .B(G122), .ZN(n453) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT107), .Z(n454) );
  XNOR2_X1 U442 ( .A(KEYINPUT102), .B(KEYINPUT12), .ZN(n462) );
  NOR2_X1 U443 ( .A1(n628), .A2(KEYINPUT65), .ZN(n410) );
  INV_X1 U444 ( .A(KEYINPUT111), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n459), .B(G478), .ZN(n556) );
  XNOR2_X1 U446 ( .A(n595), .B(KEYINPUT76), .ZN(n620) );
  AND2_X1 U447 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U448 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U449 ( .A1(n695), .A2(n605), .ZN(n594) );
  XNOR2_X1 U450 ( .A(n527), .B(n359), .ZN(n358) );
  INV_X1 U451 ( .A(KEYINPUT94), .ZN(n359) );
  BUF_X1 U452 ( .A(n538), .Z(n569) );
  BUF_X1 U453 ( .A(n755), .Z(n370) );
  XNOR2_X1 U454 ( .A(n442), .B(n352), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n363), .B(n354), .ZN(G57) );
  NAND2_X1 U456 ( .A1(n365), .A2(n364), .ZN(n363) );
  INV_X1 U457 ( .A(n738), .ZN(n364) );
  INV_X1 U458 ( .A(n711), .ZN(n400) );
  XOR2_X1 U459 ( .A(KEYINPUT110), .B(KEYINPUT6), .Z(n351) );
  XOR2_X1 U460 ( .A(n439), .B(n438), .Z(n352) );
  XNOR2_X1 U461 ( .A(n360), .B(n358), .ZN(n551) );
  XOR2_X1 U462 ( .A(n447), .B(n446), .Z(n353) );
  AND2_X1 U463 ( .A1(n711), .A2(KEYINPUT88), .ZN(n402) );
  INV_X1 U464 ( .A(n402), .ZN(n397) );
  INV_X1 U465 ( .A(KEYINPUT65), .ZN(n629) );
  XOR2_X1 U466 ( .A(KEYINPUT89), .B(KEYINPUT63), .Z(n354) );
  OR2_X2 U467 ( .A1(n585), .A2(n695), .ZN(n541) );
  XNOR2_X2 U468 ( .A(n589), .B(n351), .ZN(n585) );
  XNOR2_X2 U469 ( .A(n357), .B(n634), .ZN(n589) );
  OR2_X2 U470 ( .A1(n636), .A2(G902), .ZN(n357) );
  AND2_X1 U471 ( .A1(n734), .A2(G469), .ZN(n660) );
  AND2_X2 U472 ( .A1(n371), .A2(n633), .ZN(n734) );
  XNOR2_X2 U473 ( .A(n582), .B(KEYINPUT19), .ZN(n612) );
  XNOR2_X2 U474 ( .A(n362), .B(n361), .ZN(n481) );
  XNOR2_X2 U475 ( .A(G101), .B(KEYINPUT69), .ZN(n361) );
  XNOR2_X2 U476 ( .A(G119), .B(G113), .ZN(n362) );
  NAND2_X1 U477 ( .A1(n371), .A2(n372), .ZN(n366) );
  NOR2_X1 U478 ( .A1(n589), .A2(n400), .ZN(n590) );
  NOR2_X1 U479 ( .A1(n612), .A2(n526), .ZN(n367) );
  XNOR2_X1 U480 ( .A(n745), .B(n515), .ZN(n368) );
  XNOR2_X1 U481 ( .A(n367), .B(n527), .ZN(n369) );
  XNOR2_X1 U482 ( .A(G113), .B(G143), .ZN(n461) );
  AND2_X1 U483 ( .A1(n633), .A2(G472), .ZN(n372) );
  NAND2_X1 U484 ( .A1(n692), .A2(KEYINPUT2), .ZN(n633) );
  BUF_X1 U485 ( .A(n502), .Z(n373) );
  XOR2_X1 U486 ( .A(G140), .B(n374), .Z(n489) );
  AND2_X1 U487 ( .A1(G210), .A2(n633), .ZN(n375) );
  NAND2_X1 U488 ( .A1(n408), .A2(n407), .ZN(n391) );
  NAND2_X1 U489 ( .A1(n376), .A2(n377), .ZN(n641) );
  AND2_X1 U490 ( .A1(G475), .A2(n633), .ZN(n377) );
  AND2_X2 U491 ( .A1(n378), .A2(n409), .ZN(n379) );
  NAND2_X1 U492 ( .A1(n419), .A2(n413), .ZN(n378) );
  XNOR2_X1 U493 ( .A(n581), .B(KEYINPUT84), .ZN(n419) );
  AND2_X1 U494 ( .A1(n591), .A2(n592), .ZN(n593) );
  XNOR2_X1 U495 ( .A(n478), .B(n461), .ZN(n465) );
  XNOR2_X2 U496 ( .A(n460), .B(G131), .ZN(n478) );
  XNOR2_X1 U497 ( .A(n530), .B(n381), .ZN(n380) );
  NAND2_X1 U498 ( .A1(n623), .A2(n678), .ZN(n599) );
  XNOR2_X2 U499 ( .A(n597), .B(n598), .ZN(n623) );
  INV_X1 U500 ( .A(n611), .ZN(n386) );
  NAND2_X1 U501 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X2 U502 ( .A1(n393), .A2(n350), .ZN(n392) );
  OR2_X2 U503 ( .A1(n658), .A2(G902), .ZN(n496) );
  XNOR2_X2 U504 ( .A(n605), .B(KEYINPUT1), .ZN(n696) );
  NAND2_X1 U505 ( .A1(n401), .A2(n399), .ZN(n398) );
  NOR2_X1 U506 ( .A1(n689), .A2(n551), .ZN(n544) );
  XNOR2_X2 U507 ( .A(n496), .B(n654), .ZN(n605) );
  XNOR2_X2 U508 ( .A(n387), .B(n353), .ZN(n699) );
  NAND2_X2 U509 ( .A1(n394), .A2(n392), .ZN(n582) );
  OR2_X1 U510 ( .A1(n644), .A2(n406), .ZN(n403) );
  OR2_X1 U511 ( .A1(n368), .A2(n396), .ZN(n401) );
  OR2_X1 U512 ( .A1(n406), .A2(n397), .ZN(n396) );
  NAND2_X1 U513 ( .A1(n350), .A2(n403), .ZN(n521) );
  XNOR2_X2 U514 ( .A(KEYINPUT75), .B(n468), .ZN(n483) );
  XNOR2_X2 U515 ( .A(n479), .B(KEYINPUT4), .ZN(n513) );
  XNOR2_X2 U516 ( .A(G143), .B(G128), .ZN(n479) );
  INV_X1 U517 ( .A(n589), .ZN(n701) );
  NAND2_X1 U518 ( .A1(n375), .A2(n376), .ZN(n649) );
  NAND2_X1 U519 ( .A1(n644), .A2(n519), .ZN(n408) );
  NOR2_X1 U520 ( .A1(n411), .A2(n410), .ZN(n409) );
  NOR2_X1 U521 ( .A1(n417), .A2(n412), .ZN(n411) );
  AND2_X1 U522 ( .A1(n417), .A2(n629), .ZN(n413) );
  INV_X1 U523 ( .A(n419), .ZN(n416) );
  INV_X1 U524 ( .A(KEYINPUT74), .ZN(n418) );
  BUF_X1 U525 ( .A(n689), .Z(n720) );
  NOR2_X1 U526 ( .A1(n721), .A2(n720), .ZN(n420) );
  INV_X1 U527 ( .A(KEYINPUT46), .ZN(n609) );
  XNOR2_X1 U528 ( .A(n610), .B(n609), .ZN(n611) );
  BUF_X1 U529 ( .A(n504), .Z(n469) );
  BUF_X1 U530 ( .A(n751), .Z(n753) );
  BUF_X1 U531 ( .A(n632), .Z(n754) );
  BUF_X1 U532 ( .A(n745), .Z(n746) );
  XNOR2_X1 U533 ( .A(n421), .B(KEYINPUT14), .ZN(n422) );
  NAND2_X1 U534 ( .A1(G952), .A2(n422), .ZN(n725) );
  NOR2_X1 U535 ( .A1(n725), .A2(G953), .ZN(n524) );
  NAND2_X1 U536 ( .A1(n422), .A2(G902), .ZN(n423) );
  XNOR2_X1 U537 ( .A(n423), .B(KEYINPUT93), .ZN(n523) );
  INV_X1 U538 ( .A(n370), .ZN(n425) );
  NAND2_X1 U539 ( .A1(n523), .A2(n425), .ZN(n426) );
  NOR2_X1 U540 ( .A1(G900), .A2(n426), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n427), .B(KEYINPUT114), .ZN(n428) );
  NOR2_X1 U542 ( .A1(n524), .A2(n428), .ZN(n429) );
  XOR2_X1 U543 ( .A(KEYINPUT80), .B(n429), .Z(n592) );
  NAND2_X1 U544 ( .A1(n580), .A2(G234), .ZN(n430) );
  XNOR2_X1 U545 ( .A(n430), .B(KEYINPUT20), .ZN(n431) );
  XNOR2_X1 U546 ( .A(KEYINPUT96), .B(n431), .ZN(n444) );
  NAND2_X1 U547 ( .A1(n444), .A2(G221), .ZN(n432) );
  XNOR2_X2 U548 ( .A(G146), .B(G125), .ZN(n510) );
  XNOR2_X1 U549 ( .A(n433), .B(G140), .ZN(n434) );
  XNOR2_X1 U550 ( .A(n510), .B(n434), .ZN(n752) );
  XOR2_X1 U551 ( .A(G110), .B(G128), .Z(n436) );
  XNOR2_X1 U552 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U553 ( .A(n752), .B(n437), .ZN(n443) );
  NAND2_X1 U554 ( .A1(n755), .A2(G234), .ZN(n441) );
  NAND2_X1 U555 ( .A1(n448), .A2(G221), .ZN(n442) );
  NAND2_X1 U556 ( .A1(G217), .A2(n444), .ZN(n447) );
  XNOR2_X1 U557 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n445), .B(KEYINPUT97), .ZN(n446) );
  INV_X1 U559 ( .A(n699), .ZN(n565) );
  XNOR2_X2 U560 ( .A(G116), .B(G107), .ZN(n502) );
  XOR2_X1 U561 ( .A(n373), .B(n479), .Z(n449) );
  XNOR2_X1 U562 ( .A(n450), .B(n449), .ZN(n458) );
  XNOR2_X1 U563 ( .A(n452), .B(n451), .ZN(n456) );
  XNOR2_X1 U564 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U565 ( .A(n456), .B(n455), .Z(n457) );
  XNOR2_X1 U566 ( .A(n458), .B(n457), .ZN(n731) );
  NOR2_X1 U567 ( .A1(n731), .A2(G902), .ZN(n459) );
  XNOR2_X1 U568 ( .A(KEYINPUT13), .B(G475), .ZN(n475) );
  XNOR2_X1 U569 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U570 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U571 ( .A(n466), .B(n752), .ZN(n473) );
  INV_X1 U572 ( .A(n467), .ZN(n468) );
  NAND2_X1 U573 ( .A1(n483), .A2(G214), .ZN(n471) );
  XNOR2_X2 U574 ( .A(G122), .B(G104), .ZN(n504) );
  XNOR2_X1 U575 ( .A(n469), .B(KEYINPUT101), .ZN(n470) );
  XOR2_X1 U576 ( .A(n471), .B(n470), .Z(n472) );
  XNOR2_X1 U577 ( .A(n473), .B(n472), .ZN(n639) );
  NOR2_X1 U578 ( .A1(G902), .A2(n639), .ZN(n474) );
  NAND2_X1 U579 ( .A1(n556), .A2(n557), .ZN(n476) );
  XNOR2_X1 U580 ( .A(n476), .B(KEYINPUT108), .ZN(n676) );
  NOR2_X1 U581 ( .A1(n603), .A2(n676), .ZN(n584) );
  INV_X1 U582 ( .A(G137), .ZN(n477) );
  XNOR2_X2 U583 ( .A(n481), .B(n480), .ZN(n508) );
  XOR2_X1 U584 ( .A(n482), .B(KEYINPUT5), .Z(n485) );
  NAND2_X1 U585 ( .A1(n483), .A2(G210), .ZN(n484) );
  XNOR2_X1 U586 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n486), .B(n508), .ZN(n487) );
  XNOR2_X1 U588 ( .A(n495), .B(n487), .ZN(n636) );
  INV_X1 U589 ( .A(G472), .ZN(n634) );
  INV_X1 U590 ( .A(n348), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n584), .A2(n532), .ZN(n497) );
  XNOR2_X1 U592 ( .A(n489), .B(n488), .ZN(n491) );
  NAND2_X1 U593 ( .A1(n370), .A2(G227), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n491), .B(n490), .ZN(n493) );
  XNOR2_X2 U595 ( .A(G110), .B(KEYINPUT73), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n503), .B(KEYINPUT78), .ZN(n492) );
  XNOR2_X1 U597 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n495), .B(n494), .ZN(n658) );
  INV_X1 U599 ( .A(G469), .ZN(n654) );
  INV_X1 U600 ( .A(n696), .ZN(n567) );
  NOR2_X1 U601 ( .A1(n497), .A2(n567), .ZN(n500) );
  NAND2_X1 U602 ( .A1(n499), .A2(n498), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n516), .A2(G214), .ZN(n711) );
  NAND2_X1 U604 ( .A1(n500), .A2(n711), .ZN(n501) );
  XNOR2_X1 U605 ( .A(KEYINPUT43), .B(n501), .ZN(n520) );
  XNOR2_X1 U606 ( .A(n503), .B(n502), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n504), .B(KEYINPUT16), .ZN(n505) );
  XNOR2_X1 U608 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U609 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n510), .B(n509), .ZN(n512) );
  NAND2_X1 U611 ( .A1(n755), .A2(G224), .ZN(n511) );
  XNOR2_X1 U612 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U613 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U614 ( .A(n580), .ZN(n627) );
  NAND2_X1 U615 ( .A1(n516), .A2(G210), .ZN(n517) );
  XNOR2_X1 U616 ( .A(n517), .B(KEYINPUT92), .ZN(n518) );
  INV_X1 U617 ( .A(n518), .ZN(n519) );
  INV_X1 U618 ( .A(n521), .ZN(n596) );
  NAND2_X1 U619 ( .A1(n520), .A2(n596), .ZN(n624) );
  XNOR2_X1 U620 ( .A(n624), .B(G140), .ZN(G42) );
  INV_X1 U621 ( .A(KEYINPUT88), .ZN(n522) );
  NOR2_X1 U622 ( .A1(G898), .A2(n739), .ZN(n747) );
  AND2_X1 U623 ( .A1(n523), .A2(n747), .ZN(n525) );
  INV_X1 U624 ( .A(KEYINPUT0), .ZN(n527) );
  INV_X1 U625 ( .A(n557), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n528), .A2(n556), .ZN(n714) );
  INV_X1 U627 ( .A(n714), .ZN(n529) );
  NAND2_X1 U628 ( .A1(n529), .A2(n698), .ZN(n530) );
  INV_X1 U629 ( .A(n569), .ZN(n535) );
  NOR2_X1 U630 ( .A1(n532), .A2(n565), .ZN(n533) );
  NAND2_X1 U631 ( .A1(n533), .A2(n696), .ZN(n534) );
  NOR2_X1 U632 ( .A1(n535), .A2(n534), .ZN(n560) );
  XOR2_X1 U633 ( .A(G101), .B(n560), .Z(G3) );
  NAND2_X1 U634 ( .A1(n348), .A2(n565), .ZN(n536) );
  NOR2_X1 U635 ( .A1(n536), .A2(n696), .ZN(n537) );
  XNOR2_X1 U636 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n539) );
  XNOR2_X2 U637 ( .A(n540), .B(n539), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(G119), .ZN(G21) );
  NOR2_X1 U639 ( .A1(n541), .A2(n696), .ZN(n543) );
  XNOR2_X1 U640 ( .A(KEYINPUT112), .B(KEYINPUT33), .ZN(n542) );
  XNOR2_X1 U641 ( .A(n543), .B(n542), .ZN(n689) );
  XNOR2_X1 U642 ( .A(n544), .B(KEYINPUT34), .ZN(n547) );
  INV_X1 U643 ( .A(n556), .ZN(n545) );
  NAND2_X1 U644 ( .A1(n557), .A2(n545), .ZN(n546) );
  XNOR2_X1 U645 ( .A(n546), .B(KEYINPUT113), .ZN(n618) );
  NAND2_X1 U646 ( .A1(n547), .A2(n618), .ZN(n548) );
  XNOR2_X2 U647 ( .A(n548), .B(KEYINPUT35), .ZN(n652) );
  NAND2_X1 U648 ( .A1(n652), .A2(KEYINPUT44), .ZN(n550) );
  XNOR2_X1 U649 ( .A(n550), .B(n549), .ZN(n563) );
  INV_X1 U650 ( .A(n701), .ZN(n602) );
  NAND2_X1 U651 ( .A1(n594), .A2(n602), .ZN(n552) );
  NOR2_X1 U652 ( .A1(n551), .A2(n552), .ZN(n553) );
  XNOR2_X1 U653 ( .A(n553), .B(KEYINPUT100), .ZN(n664) );
  NOR2_X1 U654 ( .A1(n695), .A2(n602), .ZN(n554) );
  NAND2_X1 U655 ( .A1(n567), .A2(n554), .ZN(n705) );
  NOR2_X1 U656 ( .A1(n369), .A2(n705), .ZN(n555) );
  XOR2_X1 U657 ( .A(KEYINPUT31), .B(n555), .Z(n682) );
  NOR2_X1 U658 ( .A1(n664), .A2(n682), .ZN(n559) );
  NOR2_X1 U659 ( .A1(n557), .A2(n556), .ZN(n681) );
  INV_X1 U660 ( .A(n681), .ZN(n670) );
  NAND2_X1 U661 ( .A1(n670), .A2(n676), .ZN(n558) );
  XNOR2_X1 U662 ( .A(n558), .B(KEYINPUT109), .ZN(n716) );
  NOR2_X1 U663 ( .A1(n559), .A2(n716), .ZN(n561) );
  NOR2_X1 U664 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U665 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U666 ( .A(n564), .B(KEYINPUT86), .ZN(n578) );
  NAND2_X1 U667 ( .A1(n565), .A2(n602), .ZN(n566) );
  NOR2_X1 U668 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U669 ( .A1(n569), .A2(n568), .ZN(n669) );
  NAND2_X1 U670 ( .A1(n570), .A2(n669), .ZN(n574) );
  XNOR2_X1 U671 ( .A(n571), .B(KEYINPUT72), .ZN(n572) );
  NOR2_X1 U672 ( .A1(n572), .A2(KEYINPUT44), .ZN(n576) );
  NAND2_X1 U673 ( .A1(KEYINPUT72), .A2(KEYINPUT44), .ZN(n573) );
  NOR2_X1 U674 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U675 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U676 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U677 ( .A(n579), .B(KEYINPUT45), .ZN(n630) );
  NOR2_X1 U678 ( .A1(n630), .A2(n580), .ZN(n581) );
  BUF_X1 U679 ( .A(n582), .Z(n583) );
  NAND2_X1 U680 ( .A1(n584), .A2(n583), .ZN(n586) );
  NOR2_X1 U681 ( .A1(n586), .A2(n348), .ZN(n587) );
  XOR2_X1 U682 ( .A(KEYINPUT36), .B(n587), .Z(n588) );
  NOR2_X1 U683 ( .A1(n696), .A2(n588), .ZN(n685) );
  INV_X1 U684 ( .A(KEYINPUT40), .ZN(n600) );
  INV_X1 U685 ( .A(n676), .ZN(n678) );
  XOR2_X1 U686 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n598) );
  XNOR2_X1 U687 ( .A(n590), .B(KEYINPUT30), .ZN(n591) );
  XNOR2_X1 U688 ( .A(n596), .B(KEYINPUT38), .ZN(n712) );
  NAND2_X1 U689 ( .A1(n620), .A2(n712), .ZN(n597) );
  XNOR2_X1 U690 ( .A(n600), .B(n599), .ZN(n763) );
  NAND2_X1 U691 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U692 ( .A1(n714), .A2(n715), .ZN(n601) );
  XNOR2_X1 U693 ( .A(n601), .B(KEYINPUT41), .ZN(n710) );
  XNOR2_X1 U694 ( .A(n604), .B(KEYINPUT28), .ZN(n607) );
  INV_X1 U695 ( .A(n605), .ZN(n606) );
  NAND2_X1 U696 ( .A1(n607), .A2(n606), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n710), .A2(n614), .ZN(n608) );
  XNOR2_X1 U698 ( .A(n608), .B(KEYINPUT42), .ZN(n764) );
  NOR2_X1 U699 ( .A1(n763), .A2(n764), .ZN(n610) );
  BUF_X1 U700 ( .A(n612), .Z(n613) );
  NOR2_X1 U701 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U702 ( .A(n615), .B(KEYINPUT79), .ZN(n675) );
  NOR2_X1 U703 ( .A1(n716), .A2(n675), .ZN(n616) );
  XNOR2_X1 U704 ( .A(n616), .B(KEYINPUT47), .ZN(n617) );
  AND2_X1 U705 ( .A1(n521), .A2(n618), .ZN(n619) );
  NAND2_X1 U706 ( .A1(n620), .A2(n619), .ZN(n673) );
  INV_X1 U707 ( .A(KEYINPUT82), .ZN(n621) );
  XNOR2_X1 U708 ( .A(n673), .B(n621), .ZN(n622) );
  NAND2_X1 U709 ( .A1(n623), .A2(n681), .ZN(n688) );
  AND2_X1 U710 ( .A1(n688), .A2(n624), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n627), .A2(KEYINPUT2), .ZN(n628) );
  BUF_X1 U713 ( .A(n630), .Z(n631) );
  XNOR2_X1 U714 ( .A(KEYINPUT115), .B(KEYINPUT62), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n349), .B(n635), .ZN(n637) );
  OR2_X1 U716 ( .A1(n370), .A2(G952), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U718 ( .A1(n642), .A2(n738), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n643), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U720 ( .A(n368), .Z(n645) );
  XOR2_X1 U721 ( .A(KEYINPUT90), .B(KEYINPUT54), .Z(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(KEYINPUT55), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X2 U724 ( .A1(n650), .A2(n738), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U726 ( .A(n652), .Z(n653) );
  XOR2_X1 U727 ( .A(n653), .B(G122), .Z(G24) );
  XOR2_X1 U728 ( .A(KEYINPUT125), .B(KEYINPUT57), .Z(n656) );
  XNOR2_X1 U729 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n661), .A2(n738), .ZN(G54) );
  NAND2_X1 U734 ( .A1(n664), .A2(n678), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(KEYINPUT116), .ZN(n663) );
  XNOR2_X1 U736 ( .A(G104), .B(n663), .ZN(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n666) );
  NAND2_X1 U738 ( .A1(n681), .A2(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U740 ( .A(n374), .B(KEYINPUT26), .Z(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(G9) );
  XNOR2_X1 U742 ( .A(G110), .B(n669), .ZN(G12) );
  NOR2_X1 U743 ( .A1(n670), .A2(n675), .ZN(n672) );
  XNOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(G30) );
  XNOR2_X1 U746 ( .A(n673), .B(G143), .ZN(n674) );
  XNOR2_X1 U747 ( .A(KEYINPUT118), .B(n674), .ZN(G45) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U749 ( .A(G146), .B(n677), .Z(G48) );
  XOR2_X1 U750 ( .A(G113), .B(KEYINPUT119), .Z(n680) );
  NAND2_X1 U751 ( .A1(n682), .A2(n678), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(G15) );
  NAND2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n683), .B(KEYINPUT120), .ZN(n684) );
  XNOR2_X1 U755 ( .A(G116), .B(n684), .ZN(G18) );
  XNOR2_X1 U756 ( .A(G125), .B(n685), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U758 ( .A(G134), .B(KEYINPUT121), .Z(n687) );
  XNOR2_X1 U759 ( .A(n688), .B(n687), .ZN(G36) );
  NOR2_X1 U760 ( .A1(n710), .A2(n720), .ZN(n690) );
  NOR2_X1 U761 ( .A1(n690), .A2(G953), .ZN(n729) );
  NOR2_X1 U762 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n691) );
  XNOR2_X1 U763 ( .A(n692), .B(n691), .ZN(n694) );
  NAND2_X1 U764 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n693) );
  AND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n727) );
  XOR2_X1 U766 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n708) );
  NAND2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U768 ( .A(n697), .B(KEYINPUT50), .ZN(n704) );
  NOR2_X1 U769 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U770 ( .A(KEYINPUT49), .B(n700), .Z(n702) );
  NOR2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U774 ( .A(n708), .B(n707), .Z(n709) );
  NOR2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n722) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n719) );
  NOR2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U779 ( .A(KEYINPUT123), .B(n717), .Z(n718) );
  NOR2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n721) );
  NOR2_X1 U781 ( .A1(n722), .A2(n420), .ZN(n723) );
  XNOR2_X1 U782 ( .A(n723), .B(KEYINPUT52), .ZN(n724) );
  NOR2_X1 U783 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U784 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U786 ( .A(KEYINPUT53), .B(n730), .Z(G75) );
  NAND2_X1 U787 ( .A1(n734), .A2(G478), .ZN(n732) );
  XNOR2_X1 U788 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U789 ( .A1(n738), .A2(n733), .ZN(G63) );
  NAND2_X1 U790 ( .A1(n734), .A2(G217), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U792 ( .A1(n738), .A2(n737), .ZN(G66) );
  INV_X1 U793 ( .A(n631), .ZN(n740) );
  NAND2_X1 U794 ( .A1(n740), .A2(n739), .ZN(n744) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n741) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n741), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n742), .A2(G898), .ZN(n743) );
  NAND2_X1 U798 ( .A1(n744), .A2(n743), .ZN(n750) );
  XNOR2_X1 U799 ( .A(n746), .B(KEYINPUT126), .ZN(n748) );
  NOR2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U802 ( .A(n753), .B(n752), .Z(n757) );
  XNOR2_X1 U803 ( .A(n754), .B(n757), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(n370), .ZN(n761) );
  XNOR2_X1 U805 ( .A(n757), .B(G227), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U809 ( .A(KEYINPUT127), .B(n762), .Z(G72) );
  XOR2_X1 U810 ( .A(n763), .B(G131), .Z(G33) );
  XOR2_X1 U811 ( .A(G137), .B(n764), .Z(G39) );
endmodule

