

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U319 ( .A(n400), .B(KEYINPUT95), .ZN(n401) );
  INV_X1 U320 ( .A(KEYINPUT26), .ZN(n400) );
  XNOR2_X1 U321 ( .A(n413), .B(KEYINPUT37), .ZN(n414) );
  XNOR2_X1 U322 ( .A(n377), .B(n376), .ZN(n389) );
  XNOR2_X1 U323 ( .A(n365), .B(n364), .ZN(n367) );
  NOR2_X1 U324 ( .A1(n518), .A2(n538), .ZN(n522) );
  INV_X1 U325 ( .A(KEYINPUT55), .ZN(n466) );
  XNOR2_X1 U326 ( .A(n300), .B(n299), .ZN(n304) );
  XNOR2_X1 U327 ( .A(n446), .B(n445), .ZN(n496) );
  XNOR2_X1 U328 ( .A(n393), .B(n392), .ZN(n523) );
  AND2_X1 U329 ( .A1(G226GAT), .A2(G233GAT), .ZN(n287) );
  AND2_X1 U330 ( .A1(G231GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U331 ( .A(n449), .B(KEYINPUT45), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U333 ( .A(G57GAT), .B(KEYINPUT13), .Z(n440) );
  XNOR2_X1 U334 ( .A(n375), .B(KEYINPUT82), .ZN(n376) );
  XNOR2_X1 U335 ( .A(n309), .B(n288), .ZN(n310) );
  XNOR2_X1 U336 ( .A(n371), .B(n287), .ZN(n372) );
  XNOR2_X1 U337 ( .A(n311), .B(n310), .ZN(n315) );
  XNOR2_X1 U338 ( .A(n367), .B(n366), .ZN(n444) );
  XNOR2_X1 U339 ( .A(n298), .B(KEYINPUT10), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n373), .B(n372), .ZN(n379) );
  XNOR2_X1 U341 ( .A(n402), .B(n401), .ZN(n566) );
  XOR2_X1 U342 ( .A(n323), .B(n322), .Z(n531) );
  NOR2_X1 U343 ( .A1(n470), .A2(n469), .ZN(n561) );
  XOR2_X1 U344 ( .A(n392), .B(n363), .Z(n564) );
  XNOR2_X1 U345 ( .A(G183GAT), .B(KEYINPUT126), .ZN(n471) );
  XNOR2_X1 U346 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n447) );
  XNOR2_X1 U347 ( .A(n476), .B(G43GAT), .ZN(n477) );
  XNOR2_X1 U348 ( .A(n472), .B(n471), .ZN(G1350GAT) );
  XNOR2_X1 U349 ( .A(n448), .B(n447), .ZN(G1331GAT) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G99GAT), .Z(n432) );
  XOR2_X1 U351 ( .A(G162GAT), .B(G50GAT), .Z(n326) );
  XOR2_X1 U352 ( .A(n432), .B(n326), .Z(n290) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U354 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U355 ( .A(G190GAT), .B(G36GAT), .Z(n371) );
  XOR2_X1 U356 ( .A(n291), .B(n371), .Z(n300) );
  XOR2_X1 U357 ( .A(KEYINPUT71), .B(G92GAT), .Z(n293) );
  XNOR2_X1 U358 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n292) );
  XNOR2_X1 U359 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U360 ( .A(G106GAT), .B(KEYINPUT11), .Z(n295) );
  XNOR2_X1 U361 ( .A(G134GAT), .B(KEYINPUT72), .ZN(n294) );
  XNOR2_X1 U362 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U363 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U364 ( .A(G43GAT), .B(KEYINPUT7), .Z(n302) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U366 ( .A(n302), .B(n301), .ZN(n420) );
  XNOR2_X1 U367 ( .A(n420), .B(KEYINPUT73), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n560) );
  XOR2_X1 U369 ( .A(KEYINPUT36), .B(n560), .Z(n579) );
  XOR2_X1 U370 ( .A(G211GAT), .B(G78GAT), .Z(n306) );
  XNOR2_X1 U371 ( .A(n440), .B(KEYINPUT77), .ZN(n305) );
  XNOR2_X1 U372 ( .A(n306), .B(n305), .ZN(n311) );
  XOR2_X1 U373 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n308) );
  XNOR2_X1 U374 ( .A(KEYINPUT12), .B(KEYINPUT75), .ZN(n307) );
  XNOR2_X1 U375 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U376 ( .A(G183GAT), .B(G71GAT), .Z(n313) );
  XNOR2_X1 U377 ( .A(G127GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U378 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U379 ( .A(n315), .B(n314), .Z(n323) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G22GAT), .Z(n317) );
  XNOR2_X1 U381 ( .A(G8GAT), .B(KEYINPUT67), .ZN(n316) );
  XNOR2_X1 U382 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U383 ( .A(G1GAT), .B(n318), .Z(n419) );
  XOR2_X1 U384 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n320) );
  XNOR2_X1 U385 ( .A(G64GAT), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U386 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U387 ( .A(n419), .B(n321), .ZN(n322) );
  INV_X1 U388 ( .A(n531), .ZN(n576) );
  INV_X1 U389 ( .A(KEYINPUT94), .ZN(n396) );
  XOR2_X1 U390 ( .A(G197GAT), .B(KEYINPUT21), .Z(n325) );
  XNOR2_X1 U391 ( .A(G218GAT), .B(G211GAT), .ZN(n324) );
  XNOR2_X1 U392 ( .A(n325), .B(n324), .ZN(n368) );
  XOR2_X1 U393 ( .A(G204GAT), .B(n368), .Z(n328) );
  XNOR2_X1 U394 ( .A(n326), .B(G22GAT), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n333) );
  XNOR2_X1 U396 ( .A(G148GAT), .B(G106GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n329), .B(G78GAT), .ZN(n431) );
  XOR2_X1 U398 ( .A(n431), .B(KEYINPUT22), .Z(n331) );
  NAND2_X1 U399 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U400 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U401 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U402 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n335) );
  XNOR2_X1 U403 ( .A(G155GAT), .B(G141GAT), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U405 ( .A(KEYINPUT3), .B(n336), .Z(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n338) );
  XNOR2_X1 U407 ( .A(KEYINPUT86), .B(KEYINPUT84), .ZN(n337) );
  XNOR2_X1 U408 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U409 ( .A(n347), .B(n339), .ZN(n340) );
  XOR2_X1 U410 ( .A(n341), .B(n340), .Z(n399) );
  XNOR2_X1 U411 ( .A(n399), .B(KEYINPUT28), .ZN(n518) );
  XOR2_X1 U412 ( .A(KEYINPUT80), .B(G134GAT), .Z(n343) );
  XNOR2_X1 U413 ( .A(G127GAT), .B(G113GAT), .ZN(n342) );
  XNOR2_X1 U414 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U415 ( .A(KEYINPUT0), .B(n344), .ZN(n392) );
  XOR2_X1 U416 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n346) );
  XNOR2_X1 U417 ( .A(KEYINPUT88), .B(KEYINPUT91), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n348) );
  XOR2_X1 U419 ( .A(n348), .B(n347), .Z(n356) );
  XOR2_X1 U420 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n350) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U423 ( .A(G57GAT), .B(G120GAT), .Z(n352) );
  XNOR2_X1 U424 ( .A(G85GAT), .B(G148GAT), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U427 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U428 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n358) );
  NAND2_X1 U429 ( .A1(G225GAT), .A2(G233GAT), .ZN(n357) );
  XOR2_X1 U430 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U431 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U432 ( .A(G29GAT), .B(G162GAT), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U434 ( .A(G92GAT), .B(G204GAT), .ZN(n365) );
  INV_X1 U435 ( .A(G64GAT), .ZN(n364) );
  XOR2_X1 U436 ( .A(KEYINPUT70), .B(G176GAT), .Z(n366) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(n444), .Z(n370) );
  XNOR2_X1 U438 ( .A(G8GAT), .B(n368), .ZN(n369) );
  XNOR2_X1 U439 ( .A(n370), .B(n369), .ZN(n373) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n374), .B(G169GAT), .ZN(n377) );
  XNOR2_X1 U442 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n375) );
  INV_X1 U443 ( .A(n389), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n488) );
  XOR2_X1 U445 ( .A(n488), .B(KEYINPUT27), .Z(n403) );
  NAND2_X1 U446 ( .A1(n564), .A2(n403), .ZN(n538) );
  XNOR2_X1 U447 ( .A(KEYINPUT93), .B(n522), .ZN(n394) );
  XOR2_X1 U448 ( .A(KEYINPUT83), .B(KEYINPUT64), .Z(n381) );
  XNOR2_X1 U449 ( .A(G99GAT), .B(G15GAT), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U451 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XOR2_X1 U452 ( .A(n382), .B(n439), .Z(n384) );
  XNOR2_X1 U453 ( .A(G43GAT), .B(G190GAT), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U455 ( .A(KEYINPUT81), .B(G176GAT), .Z(n386) );
  NAND2_X1 U456 ( .A1(G227GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U457 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U458 ( .A(n388), .B(n387), .Z(n391) );
  XOR2_X1 U459 ( .A(n389), .B(KEYINPUT20), .Z(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n393) );
  NOR2_X1 U461 ( .A1(n394), .A2(n523), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n410) );
  INV_X1 U463 ( .A(n523), .ZN(n470) );
  NOR2_X1 U464 ( .A1(n470), .A2(n488), .ZN(n397) );
  NOR2_X1 U465 ( .A1(n399), .A2(n397), .ZN(n398) );
  XOR2_X1 U466 ( .A(KEYINPUT25), .B(n398), .Z(n406) );
  INV_X1 U467 ( .A(n399), .ZN(n464) );
  NOR2_X1 U468 ( .A1(n464), .A2(n523), .ZN(n402) );
  AND2_X1 U469 ( .A1(n566), .A2(n403), .ZN(n404) );
  XNOR2_X1 U470 ( .A(KEYINPUT96), .B(n404), .ZN(n405) );
  NOR2_X1 U471 ( .A1(n406), .A2(n405), .ZN(n407) );
  NOR2_X1 U472 ( .A1(n407), .A2(n564), .ZN(n408) );
  XNOR2_X1 U473 ( .A(KEYINPUT97), .B(n408), .ZN(n409) );
  NAND2_X1 U474 ( .A1(n410), .A2(n409), .ZN(n481) );
  NAND2_X1 U475 ( .A1(n576), .A2(n481), .ZN(n411) );
  XOR2_X1 U476 ( .A(KEYINPUT103), .B(n411), .Z(n412) );
  NOR2_X1 U477 ( .A1(n579), .A2(n412), .ZN(n415) );
  XOR2_X1 U478 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n413) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n510) );
  XOR2_X1 U480 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n417) );
  XNOR2_X1 U481 ( .A(G113GAT), .B(G169GAT), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n430) );
  XOR2_X1 U484 ( .A(G197GAT), .B(G50GAT), .Z(n422) );
  XNOR2_X1 U485 ( .A(n420), .B(G36GAT), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U487 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n424) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U490 ( .A(n426), .B(n425), .Z(n428) );
  XNOR2_X1 U491 ( .A(G141GAT), .B(KEYINPUT65), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U493 ( .A(n430), .B(n429), .Z(n568) );
  INV_X1 U494 ( .A(n568), .ZN(n552) );
  XOR2_X1 U495 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT69), .B(KEYINPUT31), .Z(n436) );
  XNOR2_X1 U499 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U501 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n572) );
  NAND2_X1 U505 ( .A1(n552), .A2(n572), .ZN(n484) );
  NOR2_X1 U506 ( .A1(n510), .A2(n484), .ZN(n446) );
  XNOR2_X1 U507 ( .A(KEYINPUT38), .B(KEYINPUT106), .ZN(n445) );
  NAND2_X1 U508 ( .A1(n496), .A2(n518), .ZN(n448) );
  INV_X1 U509 ( .A(KEYINPUT54), .ZN(n463) );
  NOR2_X1 U510 ( .A1(n576), .A2(n579), .ZN(n451) );
  INV_X1 U511 ( .A(KEYINPUT115), .ZN(n449) );
  NAND2_X1 U512 ( .A1(n452), .A2(n572), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(KEYINPUT116), .ZN(n454) );
  NOR2_X1 U514 ( .A1(n454), .A2(n552), .ZN(n460) );
  INV_X1 U515 ( .A(n560), .ZN(n550) );
  NAND2_X1 U516 ( .A1(n550), .A2(n576), .ZN(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT41), .B(n572), .Z(n541) );
  INV_X1 U518 ( .A(n541), .ZN(n557) );
  NAND2_X1 U519 ( .A1(n552), .A2(n557), .ZN(n455) );
  XOR2_X1 U520 ( .A(KEYINPUT46), .B(n455), .Z(n456) );
  NOR2_X1 U521 ( .A1(n457), .A2(n456), .ZN(n458) );
  XOR2_X1 U522 ( .A(KEYINPUT47), .B(n458), .Z(n459) );
  NOR2_X1 U523 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U524 ( .A(KEYINPUT48), .B(n461), .ZN(n537) );
  NOR2_X1 U525 ( .A1(n488), .A2(n537), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n565) );
  OR2_X1 U527 ( .A1(n564), .A2(n399), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n565), .A2(n465), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT123), .B(n468), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n531), .A2(n561), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n496), .A2(n564), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(G29GAT), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  NAND2_X1 U536 ( .A1(n496), .A2(n523), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n476) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  NAND2_X1 U539 ( .A1(n531), .A2(n550), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT79), .ZN(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT16), .B(n480), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(KEYINPUT98), .ZN(n499) );
  NOR2_X1 U544 ( .A1(n499), .A2(n484), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT99), .B(n485), .Z(n493) );
  NAND2_X1 U546 ( .A1(n564), .A2(n493), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n486), .B(KEYINPUT34), .ZN(n487) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  INV_X1 U549 ( .A(n488), .ZN(n513) );
  NAND2_X1 U550 ( .A1(n493), .A2(n513), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT100), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U554 ( .A1(n493), .A2(n523), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  XOR2_X1 U556 ( .A(G22GAT), .B(KEYINPUT101), .Z(n495) );
  NAND2_X1 U557 ( .A1(n493), .A2(n518), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(G1327GAT) );
  NAND2_X1 U559 ( .A1(n496), .A2(n513), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n501) );
  NAND2_X1 U562 ( .A1(n568), .A2(n557), .ZN(n498) );
  XOR2_X1 U563 ( .A(KEYINPUT109), .B(n498), .Z(n509) );
  NOR2_X1 U564 ( .A1(n499), .A2(n509), .ZN(n506) );
  NAND2_X1 U565 ( .A1(n506), .A2(n564), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n506), .A2(n513), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n502), .B(KEYINPUT110), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(n503), .ZN(G1333GAT) );
  XOR2_X1 U570 ( .A(G71GAT), .B(KEYINPUT111), .Z(n505) );
  NAND2_X1 U571 ( .A1(n506), .A2(n523), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U574 ( .A1(n506), .A2(n518), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n564), .A2(n519), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(KEYINPUT112), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  XOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT113), .Z(n515) );
  NAND2_X1 U581 ( .A1(n519), .A2(n513), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n523), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n516), .B(KEYINPUT114), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n517), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(G113GAT), .B(KEYINPUT117), .Z(n526) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n537), .A2(n524), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n534), .A2(n552), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U595 ( .A1(n534), .A2(n557), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n530) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT118), .Z(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n531), .A2(n534), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n560), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n539), .A2(n566), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n568), .A2(n549), .ZN(n540) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n541), .A2(n549), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n543) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(KEYINPUT52), .B(n544), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n576), .A2(n549), .ZN(n547) );
  XOR2_X1 U616 ( .A(KEYINPUT122), .B(n547), .Z(n548) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n561), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n555) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(n556), .Z(n559) );
  NAND2_X1 U626 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n578) );
  NOR2_X1 U633 ( .A1(n568), .A2(n578), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n578), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

