//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n187));
  INV_X1    g001(.A(G472), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  AOI21_X1  g005(.A(G131), .B1(new_n190), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(G137), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT67), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  OAI211_X1 g019(.A(G128), .B(new_n202), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n207), .B(new_n208), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n197), .A2(new_n198), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n200), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT68), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n200), .A2(new_n211), .A3(new_n219), .A4(new_n216), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n207), .A2(new_n208), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n191), .A2(new_n194), .A3(new_n198), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n215), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT30), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n218), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n215), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n222), .B(KEYINPUT64), .C1(new_n223), .C2(new_n224), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n191), .A2(new_n194), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n199), .B1(new_n237), .B2(new_n192), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(KEYINPUT65), .A3(new_n210), .A4(new_n206), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n206), .A2(new_n210), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n213), .A2(new_n215), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n236), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n229), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G116), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n249), .A3(G119), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n254), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n250), .A3(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n231), .A2(new_n245), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n228), .A2(new_n258), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n218), .A2(new_n260), .A3(new_n220), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT29), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT28), .B1(new_n260), .B2(new_n217), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n244), .A2(new_n258), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n261), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n267), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n218), .A2(new_n220), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n258), .B1(new_n276), .B2(new_n228), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n261), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n270), .B(KEYINPUT73), .Z(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT29), .A4(new_n267), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n188), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT70), .B1(new_n273), .B2(new_n267), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n261), .B2(new_n271), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n285), .B(new_n268), .C1(new_n287), .C2(new_n270), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n261), .A2(new_n267), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n259), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n290), .B2(new_n259), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n290), .A2(new_n259), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n293), .A3(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n289), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G472), .A2(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n283), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n304));
  INV_X1    g118(.A(new_n301), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n295), .B1(new_n293), .B2(new_n292), .ZN(new_n306));
  INV_X1    g120(.A(new_n299), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n308), .B2(new_n289), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n300), .A2(new_n301), .ZN(new_n312));
  INV_X1    g126(.A(new_n310), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT72), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n303), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(G234), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n204), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n251), .B2(G128), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n251), .A2(G128), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT76), .A4(new_n332), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(G110), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT74), .B1(new_n209), .B2(G119), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n251), .A3(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n209), .A2(G119), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT24), .B(G110), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(KEYINPUT75), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n328), .A2(new_n337), .A3(new_n345), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n320), .A2(new_n322), .A3(new_n204), .ZN(new_n350));
  INV_X1    g164(.A(G110), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n330), .A2(new_n331), .A3(new_n351), .A4(new_n332), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n342), .A2(new_n344), .B1(new_n352), .B2(KEYINPUT77), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(KEYINPUT77), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n327), .B(new_n350), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G137), .ZN(new_n356));
  INV_X1    g170(.A(G953), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(G221), .A3(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n349), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n349), .B2(new_n355), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT25), .B1(new_n362), .B2(new_n317), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n355), .ZN(new_n364));
  INV_X1    g178(.A(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n349), .A2(new_n355), .A3(new_n359), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n317), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n318), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n318), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT78), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n374));
  INV_X1    g188(.A(new_n318), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n366), .A2(new_n317), .A3(new_n367), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n378), .B2(new_n368), .ZN(new_n379));
  INV_X1    g193(.A(new_n372), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n374), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n373), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n187), .B1(new_n315), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n282), .B1(new_n309), .B2(KEYINPUT32), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT72), .B1(new_n312), .B2(new_n313), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n304), .B(new_n310), .C1(new_n300), .C2(new_n301), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n382), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(KEYINPUT79), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT9), .B(G234), .ZN(new_n390));
  OAI21_X1  g204(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G469), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(new_n317), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(G107), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(KEYINPUT81), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  INV_X1    g215(.A(new_n398), .ZN(new_n402));
  NOR2_X1   g216(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n403));
  OAI22_X1  g217(.A1(new_n402), .A2(new_n403), .B1(new_n396), .B2(G107), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n396), .A3(G107), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n400), .A2(new_n401), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G107), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n397), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n206), .A2(new_n210), .A3(new_n410), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n411), .A2(new_n241), .B1(new_n413), .B2(new_n407), .ZN(new_n414));
  INV_X1    g228(.A(new_n234), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n395), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n211), .B1(new_n407), .B2(new_n410), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n398), .A2(G104), .A3(new_n408), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT81), .B1(new_n408), .B2(G104), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n406), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n423), .A2(new_n398), .B1(G104), .B2(new_n408), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n420), .A2(new_n424), .A3(G101), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(new_n412), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT12), .B(new_n234), .C1(new_n417), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G101), .B1(new_n420), .B2(new_n424), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n407), .A2(new_n429), .A3(KEYINPUT4), .ZN(new_n430));
  INV_X1    g244(.A(new_n225), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(G101), .C1(new_n420), .C2(new_n424), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n413), .A2(KEYINPUT10), .A3(new_n407), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n425), .B2(new_n412), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n434), .A2(new_n415), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n357), .A2(G227), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n440), .B(new_n441), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n435), .A2(new_n437), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n434), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n234), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n439), .A2(new_n442), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n394), .B1(new_n448), .B2(G469), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n415), .B1(new_n445), .B2(new_n434), .ZN(new_n450));
  AND4_X1   g264(.A1(new_n415), .A2(new_n434), .A3(new_n435), .A4(new_n437), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n442), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n443), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n428), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT83), .B1(new_n438), .B2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n393), .A3(new_n317), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n392), .B1(new_n449), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G113), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n396), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT19), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT19), .B1(new_n320), .B2(new_n322), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n204), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(KEYINPUT85), .A2(G143), .ZN(new_n464));
  NOR2_X1   g278(.A1(KEYINPUT85), .A2(G143), .ZN(new_n465));
  OAI211_X1 g279(.A(G214), .B(new_n263), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G237), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n357), .A3(G214), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT85), .A2(G143), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n466), .A2(new_n196), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n196), .B1(new_n466), .B2(new_n470), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n327), .B(new_n463), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(KEYINPUT86), .A3(new_n470), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT18), .A2(G131), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT86), .A4(new_n475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n320), .A2(new_n322), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G146), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n350), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n460), .B1(new_n473), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT17), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n470), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT17), .A3(G131), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n327), .A3(new_n326), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n460), .B(new_n482), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n490), .A2(KEYINPUT87), .A3(new_n491), .A4(new_n492), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n487), .A2(new_n327), .A3(new_n326), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n486), .A2(G131), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n466), .A2(new_n196), .A3(new_n470), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n474), .A2(new_n476), .B1(new_n350), .B2(new_n480), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n497), .A2(new_n501), .B1(new_n478), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n483), .B1(new_n503), .B2(new_n460), .ZN(new_n504));
  INV_X1    g318(.A(new_n492), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT20), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n495), .A2(new_n496), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n489), .ZN(new_n508));
  INV_X1    g322(.A(new_n327), .ZN(new_n509));
  AOI21_X1  g323(.A(G146), .B1(new_n323), .B2(new_n324), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n501), .A2(new_n511), .A3(new_n487), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n460), .B1(new_n512), .B2(new_n482), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n317), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G475), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n201), .A2(G128), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n209), .A2(KEYINPUT88), .A3(G143), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT88), .B1(new_n209), .B2(G143), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G134), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n190), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT14), .A4(G122), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n247), .A2(new_n249), .A3(G122), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n246), .A2(G122), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(G107), .B(new_n524), .C1(new_n527), .C2(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n408), .A3(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n518), .B2(new_n519), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n532), .A3(G134), .ZN(new_n533));
  OAI221_X1 g347(.A(new_n517), .B1(new_n531), .B2(new_n190), .C1(new_n518), .C2(new_n519), .ZN(new_n534));
  INV_X1    g348(.A(new_n529), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n408), .B1(new_n525), .B2(new_n526), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n533), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n390), .A2(new_n316), .A3(G953), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n530), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n530), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n317), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G478), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT89), .B(new_n317), .C1(new_n539), .C2(new_n540), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n357), .A2(G952), .ZN(new_n548));
  NAND2_X1  g362(.A1(G234), .A2(G237), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(G902), .A3(G953), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT21), .B(G898), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n541), .A2(new_n545), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n547), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n516), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G214), .B1(G237), .B2(G902), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT84), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n430), .A2(new_n258), .A3(new_n433), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT5), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n251), .A3(G116), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(G113), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n253), .B2(new_n565), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n568), .A2(new_n257), .A3(new_n407), .A4(new_n410), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G122), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n569), .A3(new_n571), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(KEYINPUT6), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n241), .A2(new_n321), .ZN(new_n576));
  INV_X1    g390(.A(G224), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(G953), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n225), .A2(G125), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n576), .B2(new_n580), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT6), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n570), .A2(new_n584), .A3(new_n572), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n575), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  OAI22_X1  g400(.A1(new_n581), .A2(new_n582), .B1(KEYINPUT7), .B2(new_n578), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n571), .B(KEYINPUT8), .ZN(new_n588));
  INV_X1    g402(.A(new_n569), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n568), .A2(new_n257), .B1(new_n407), .B2(new_n410), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n576), .A2(new_n580), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n579), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n587), .A2(new_n591), .A3(new_n574), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n317), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n563), .B1(new_n586), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n595), .A2(new_n317), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n575), .A2(new_n583), .A3(new_n585), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n562), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n561), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n458), .A2(new_n559), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n383), .A2(new_n389), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n300), .A2(new_n317), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n605), .A2(G472), .B1(new_n301), .B2(new_n300), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n449), .A2(new_n457), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n391), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n382), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n530), .A2(new_n537), .ZN(new_n611));
  INV_X1    g425(.A(new_n538), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n530), .A2(new_n537), .A3(new_n538), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT33), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n544), .B1(new_n619), .B2(new_n317), .ZN(new_n620));
  AOI21_X1  g434(.A(G478), .B1(new_n543), .B2(new_n546), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT90), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n621), .ZN(new_n623));
  INV_X1    g437(.A(new_n618), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n617), .B1(new_n613), .B2(new_n614), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n317), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G478), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT90), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n516), .ZN(new_n631));
  INV_X1    g445(.A(new_n601), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n631), .A2(new_n632), .A3(new_n555), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n610), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n547), .A2(new_n557), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n555), .B(KEYINPUT91), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n506), .A2(new_n493), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n637), .A2(new_n515), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT92), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n639), .A2(new_n515), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT92), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n637), .A4(new_n638), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(new_n644), .A3(new_n601), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT93), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(new_n644), .A3(KEYINPUT93), .A4(new_n601), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n610), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n365), .A2(KEYINPUT36), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n364), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n349), .A2(new_n355), .A3(new_n653), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n371), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT94), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT94), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(new_n659), .A3(new_n371), .A4(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n370), .A2(new_n662), .A3(KEYINPUT95), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT95), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n379), .B2(new_n661), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT96), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT96), .B1(new_n663), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n606), .A2(new_n668), .A3(new_n602), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  OR2_X1    g485(.A1(new_n552), .A2(G900), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n550), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n642), .A2(new_n637), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT96), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT95), .B1(new_n370), .B2(new_n662), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n379), .A2(new_n661), .A3(new_n664), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT96), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n458), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n632), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n387), .A2(new_n675), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XNOR2_X1  g498(.A(new_n673), .B(KEYINPUT39), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n458), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n686), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n598), .A2(new_n599), .A3(new_n562), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n562), .B1(new_n598), .B2(new_n599), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n677), .A2(new_n678), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n561), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n516), .A2(new_n637), .A3(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n689), .A2(new_n692), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n311), .A2(new_n314), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT97), .ZN(new_n704));
  INV_X1    g518(.A(new_n278), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n704), .B1(new_n705), .B2(new_n267), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n278), .A2(KEYINPUT97), .A3(new_n268), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n298), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n188), .B1(new_n708), .B2(new_n317), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n309), .B2(KEYINPUT32), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n702), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n201), .ZN(G45));
  NAND3_X1  g529(.A1(new_n630), .A2(new_n516), .A3(new_n673), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n387), .A2(new_n682), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  NAND2_X1  g533(.A1(new_n456), .A2(new_n317), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(KEYINPUT100), .A3(new_n457), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n723), .A3(G469), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n392), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(new_n388), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n387), .A2(new_n726), .A3(new_n633), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT101), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n387), .A2(new_n726), .A3(new_n729), .A4(new_n633), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND3_X1  g547(.A1(new_n387), .A2(new_n649), .A3(new_n726), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  AND2_X1   g549(.A1(new_n668), .A2(new_n559), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n722), .A2(new_n724), .ZN(new_n737));
  AND4_X1   g551(.A1(KEYINPUT102), .A2(new_n737), .A3(new_n391), .A4(new_n601), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT102), .B1(new_n725), .B2(new_n601), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n387), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  OR3_X1    g556(.A1(new_n700), .A2(new_n695), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n742), .B1(new_n700), .B2(new_n695), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n188), .B1(new_n300), .B2(new_n317), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n370), .A2(new_n372), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n280), .B1(new_n705), .B2(new_n286), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n268), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n296), .A2(new_n292), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n305), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n746), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n745), .A2(new_n638), .A3(new_n725), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NOR4_X1   g568(.A1(new_n716), .A2(new_n746), .A3(new_n697), .A4(new_n751), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n738), .B2(new_n739), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  OR2_X1    g571(.A1(new_n309), .A2(KEYINPUT32), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n747), .B1(new_n758), .B2(new_n384), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n693), .A2(new_n694), .A3(new_n561), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n608), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n717), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n609), .A2(new_n760), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n315), .A2(new_n716), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n765), .B2(KEYINPUT42), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR3_X1   g581(.A1(new_n761), .A2(new_n608), .A3(new_n382), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n387), .A2(new_n675), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n516), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n630), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT43), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n516), .A2(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n516), .A2(KEYINPUT106), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n630), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n772), .B2(KEYINPUT105), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n774), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n605), .A2(G472), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n312), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n698), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT107), .B1(new_n782), .B2(new_n698), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n761), .B1(new_n787), .B2(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n444), .A2(new_n447), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n451), .B1(new_n427), .B2(new_n416), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n790), .B2(new_n443), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n448), .A2(KEYINPUT45), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(G469), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT104), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT104), .A4(G469), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n394), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n457), .B1(new_n799), .B2(KEYINPUT46), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n391), .B(new_n685), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n802), .B1(new_n786), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n788), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n391), .B1(new_n800), .B2(new_n801), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(KEYINPUT47), .B(new_n391), .C1(new_n800), .C2(new_n801), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n717), .A2(new_n382), .A3(new_n760), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n387), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n807), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(KEYINPUT108), .B(new_n814), .C1(new_n810), .C2(new_n811), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n319), .ZN(G42));
  NOR2_X1   g633(.A1(G952), .A2(G953), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT119), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n780), .A2(new_n551), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n725), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n761), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n759), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT48), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n826), .A2(KEYINPUT118), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n823), .A2(new_n752), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n830), .B1(new_n739), .B2(new_n738), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n713), .A2(new_n712), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n824), .A2(new_n382), .A3(new_n550), .A4(new_n761), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n831), .B(new_n548), .C1(new_n631), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n828), .B(new_n835), .C1(new_n826), .C2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n830), .A2(KEYINPUT116), .A3(new_n760), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n829), .B2(new_n761), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n391), .B1(new_n722), .B2(new_n724), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n838), .B(new_n840), .C1(new_n812), .C2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n696), .A2(new_n725), .A3(new_n561), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT50), .B1(new_n829), .B2(new_n843), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n829), .A2(KEYINPUT50), .A3(new_n843), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n630), .A2(new_n516), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n832), .A2(new_n833), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n746), .A2(new_n697), .A3(new_n751), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n823), .A2(new_n849), .A3(new_n825), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n848), .A2(KEYINPUT117), .A3(new_n850), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n846), .A2(new_n851), .ZN(new_n856));
  OAI221_X1 g670(.A(new_n837), .B1(new_n846), .B2(new_n855), .C1(new_n856), .C2(KEYINPUT51), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n699), .B(new_n638), .C1(new_n693), .C2(new_n694), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n637), .A2(new_n507), .A3(new_n515), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n609), .A2(new_n781), .A3(new_n860), .A4(new_n312), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT110), .B1(new_n669), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n669), .A2(new_n861), .A3(KEYINPUT110), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n631), .A2(new_n858), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n863), .A2(new_n864), .B1(new_n610), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  INV_X1    g681(.A(new_n673), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n514), .B2(G475), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n639), .A2(new_n547), .A3(new_n557), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT111), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n482), .B1(new_n485), .B2(new_n488), .ZN(new_n873));
  INV_X1    g687(.A(new_n460), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(G902), .B1(new_n875), .B2(new_n489), .ZN(new_n876));
  INV_X1    g690(.A(G475), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n673), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n493), .B2(new_n506), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(KEYINPUT111), .A3(new_n557), .A4(new_n547), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n760), .A2(new_n872), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n760), .A2(new_n880), .A3(KEYINPUT112), .A4(new_n872), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n681), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n387), .A2(new_n885), .B1(new_n755), .B2(new_n762), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n867), .B1(new_n886), .B2(new_n769), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n387), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n849), .A2(new_n717), .A3(new_n762), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n867), .A2(new_n769), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n603), .B(new_n866), .C1(new_n887), .C2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n740), .A2(new_n734), .A3(new_n753), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n731), .A3(new_n766), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT114), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n731), .A3(new_n766), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT114), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n383), .A2(new_n389), .A3(new_n602), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n610), .A2(new_n865), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n669), .A2(new_n861), .A3(KEYINPUT110), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n862), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n681), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n870), .B(KEYINPUT111), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT112), .B1(new_n903), .B2(new_n760), .ZN(new_n904));
  INV_X1    g718(.A(new_n884), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n889), .B1(new_n906), .B2(new_n315), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n315), .A2(new_n674), .A3(new_n764), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT113), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n886), .A2(new_n867), .A3(new_n769), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n895), .A2(new_n896), .A3(new_n901), .A4(new_n911), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n608), .A2(new_n379), .A3(new_n661), .A4(new_n868), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n711), .A2(new_n745), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n756), .A3(new_n683), .A4(new_n718), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT52), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n894), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n756), .A2(new_n683), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n919), .B2(KEYINPUT52), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n740), .A2(new_n734), .A3(new_n753), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n730), .B2(new_n728), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n901), .A3(new_n911), .A4(new_n766), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n916), .B1(new_n924), .B2(KEYINPUT114), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n925), .B2(new_n912), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n923), .B2(new_n766), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n893), .A2(KEYINPUT115), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n919), .B2(KEYINPUT52), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n901), .A2(new_n911), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n917), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n927), .B1(KEYINPUT54), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n821), .B1(new_n857), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n777), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n747), .A2(new_n392), .A3(new_n561), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT49), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n737), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT109), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n737), .A2(new_n942), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n944), .A2(new_n832), .A3(new_n696), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n939), .A2(new_n946), .ZN(G75));
  NOR2_X1   g761(.A1(new_n357), .A2(G952), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT120), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n937), .A2(G902), .ZN(new_n952));
  INV_X1    g766(.A(G210), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n575), .A2(new_n585), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(new_n583), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT55), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n951), .B(new_n957), .C1(new_n952), .C2(new_n953), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n959), .B2(new_n960), .ZN(G51));
  XNOR2_X1  g775(.A(new_n394), .B(KEYINPUT57), .ZN(new_n962));
  INV_X1    g776(.A(new_n934), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n895), .A2(new_n930), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n893), .A2(KEYINPUT115), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n917), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n926), .A2(new_n966), .A3(KEYINPUT54), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT54), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n929), .B2(new_n936), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n456), .ZN(new_n971));
  INV_X1    g785(.A(new_n952), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n797), .A3(new_n798), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n948), .B1(new_n971), .B2(new_n973), .ZN(G54));
  NAND2_X1  g788(.A1(KEYINPUT58), .A2(G475), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n504), .B1(new_n952), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n948), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n952), .A2(new_n504), .A3(new_n975), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G60));
  NAND2_X1  g794(.A1(G478), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT59), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n619), .B1(new_n938), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n619), .B(new_n983), .C1(new_n967), .C2(new_n969), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n949), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(G63));
  AND2_X1   g801(.A1(new_n655), .A2(new_n656), .ZN(new_n988));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n988), .B(new_n991), .C1(new_n926), .C2(new_n966), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT122), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT122), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n937), .A2(new_n994), .A3(new_n988), .A4(new_n991), .ZN(new_n995));
  INV_X1    g809(.A(new_n362), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n928), .A2(new_n918), .B1(new_n935), .B2(new_n917), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n990), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n993), .A2(new_n995), .A3(new_n949), .A4(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n998), .A2(KEYINPUT61), .A3(new_n949), .A4(new_n992), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n554), .B2(new_n577), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n923), .A2(new_n901), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n955), .B1(G898), .B2(new_n357), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G69));
  NAND2_X1  g822(.A1(new_n231), .A2(new_n245), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n461), .A2(new_n462), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n383), .A2(new_n389), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n761), .B(new_n691), .C1(new_n631), .C2(new_n859), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT124), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT124), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n805), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1018), .A2(new_n818), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n756), .A2(new_n683), .A3(new_n718), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n714), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT62), .ZN(new_n1022));
  OAI21_X1  g836(.A(KEYINPUT123), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT123), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1024), .B(KEYINPUT62), .C1(new_n714), .C2(new_n1020), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n714), .A2(new_n1020), .A3(KEYINPUT62), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1019), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1011), .B1(new_n1029), .B2(new_n357), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n816), .A2(new_n817), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1020), .B1(new_n788), .B2(new_n804), .ZN(new_n1032));
  INV_X1    g846(.A(new_n802), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1033), .A2(new_n745), .A3(new_n759), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n1034), .A2(new_n766), .A3(new_n769), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1031), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1036), .A2(G953), .ZN(new_n1037));
  NAND2_X1  g851(.A1(G900), .A2(G953), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1011), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(KEYINPUT125), .B1(new_n1030), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g855(.A(new_n1011), .B(new_n1038), .C1(new_n1036), .C2(G953), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT125), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1018), .A2(new_n818), .A3(new_n1027), .ZN(new_n1044));
  AOI21_X1  g858(.A(G953), .B1(new_n1044), .B2(new_n1026), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1042), .B(new_n1043), .C1(new_n1045), .C2(new_n1011), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n357), .B1(G227), .B2(G900), .ZN(new_n1047));
  AND3_X1   g861(.A1(new_n1041), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1047), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1048), .A2(new_n1049), .ZN(G72));
  NAND2_X1  g864(.A1(G472), .A2(G902), .ZN(new_n1051));
  XOR2_X1   g865(.A(new_n1051), .B(KEYINPUT63), .Z(new_n1052));
  INV_X1    g866(.A(new_n1005), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1052), .B1(new_n1029), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1054), .A2(new_n267), .A3(new_n262), .ZN(new_n1055));
  INV_X1    g869(.A(new_n262), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n298), .B1(new_n1056), .B2(new_n267), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(new_n1052), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT127), .Z(new_n1059));
  OAI21_X1  g873(.A(new_n1059), .B1(new_n921), .B2(new_n926), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g875(.A(KEYINPUT126), .ZN(new_n1062));
  OR2_X1    g876(.A1(new_n1036), .A2(new_n1053), .ZN(new_n1063));
  AOI211_X1 g877(.A(new_n267), .B(new_n262), .C1(new_n1063), .C2(new_n1052), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1062), .B1(new_n1064), .B2(new_n948), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1063), .A2(new_n1052), .ZN(new_n1066));
  NAND4_X1  g880(.A1(new_n1066), .A2(new_n261), .A3(new_n268), .A4(new_n259), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n1067), .A2(KEYINPUT126), .A3(new_n977), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1061), .B1(new_n1065), .B2(new_n1068), .ZN(G57));
endmodule


