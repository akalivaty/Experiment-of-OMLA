//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR3_X1   g0013(.A1(new_n212), .A2(new_n213), .A3(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G116), .A2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n222), .B(new_n227), .C1(G97), .C2(G257), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(G1), .B2(G20), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT1), .Z(new_n230));
  AOI211_X1 g0030(.A(new_n216), .B(new_n230), .C1(new_n211), .C2(new_n215), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XOR2_X1   g0047(.A(KEYINPUT8), .B(G58), .Z(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n248), .A2(new_n250), .B1(G20), .B2(new_n203), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(new_n206), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n202), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n257), .B1(G1), .B2(new_n213), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n259), .B(new_n264), .C1(new_n202), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G223), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G222), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n206), .B1(G33), .B2(G41), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n273), .B(new_n274), .C1(G77), .C2(new_n269), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n275), .B(new_n279), .C1(new_n224), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  INV_X1    g0083(.A(G190), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n266), .A2(new_n267), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n268), .A2(new_n283), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT10), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n282), .A2(G179), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n266), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n279), .B1(new_n281), .B2(new_n219), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT65), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G238), .A2(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n269), .B(new_n296), .C1(new_n233), .C2(G1698), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n274), .C1(G107), .C2(new_n269), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT15), .B(G87), .Z(new_n303));
  AOI22_X1  g0103(.A1(new_n253), .A2(new_n248), .B1(new_n303), .B2(new_n250), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n213), .B2(new_n218), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n258), .B1(new_n218), .B2(new_n263), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n265), .A2(new_n218), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n302), .B(new_n309), .C1(G169), .C2(new_n300), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n288), .A2(new_n292), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n213), .A2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n250), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n313), .B1(new_n254), .B2(new_n202), .C1(new_n314), .C2(new_n218), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT68), .B(KEYINPUT11), .Z(new_n316));
  AND3_X1   g0116(.A1(new_n315), .A2(new_n258), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n315), .B2(new_n258), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n261), .A2(new_n312), .A3(KEYINPUT12), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n225), .B2(new_n265), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT12), .B1(new_n261), .B2(new_n312), .ZN(new_n321));
  NOR4_X1   g0121(.A1(new_n317), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n233), .A2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G226), .B2(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n325), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n278), .B1(new_n332), .B2(new_n274), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n226), .B2(new_n281), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n324), .B1(new_n337), .B2(G169), .ZN(new_n338));
  AOI211_X1 g0138(.A(KEYINPUT14), .B(new_n290), .C1(new_n335), .C2(new_n336), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n337), .A2(new_n301), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n323), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n337), .A2(G200), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n322), .C1(new_n284), .C2(new_n337), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n300), .A2(G190), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n299), .A2(G200), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT72), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT16), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT69), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT69), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n269), .B2(G20), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n225), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G58), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n225), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n201), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n253), .A2(G159), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n353), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT7), .B1(new_n269), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n331), .A2(new_n358), .A3(new_n213), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(G68), .ZN(new_n370));
  INV_X1    g0170(.A(new_n366), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n258), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n224), .A2(G1698), .ZN(new_n374));
  OR2_X1    g0174(.A1(G223), .A2(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n269), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n278), .B1(new_n378), .B2(new_n274), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n280), .A2(G232), .A3(new_n276), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G200), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n265), .A2(new_n248), .ZN(new_n383));
  INV_X1    g0183(.A(new_n248), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n262), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT70), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(KEYINPUT70), .A3(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(G190), .A3(new_n380), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n373), .A2(new_n382), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n352), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n392), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(new_n393), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(KEYINPUT72), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n373), .A2(new_n390), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n373), .A2(new_n390), .A3(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n290), .B1(new_n379), .B2(new_n380), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n301), .B2(new_n381), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT18), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n381), .A2(new_n301), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n406), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n410), .B(new_n412), .C1(new_n403), .C2(new_n404), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n396), .B(new_n400), .C1(new_n409), .C2(new_n413), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n311), .A2(new_n345), .A3(new_n351), .A4(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G20), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT23), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n269), .A2(new_n213), .A3(G87), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT22), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT22), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n269), .A2(new_n422), .A3(new_n213), .A4(G87), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT24), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n250), .A2(G116), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n258), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n212), .A2(G33), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n257), .A2(new_n262), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G107), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n418), .A2(G1), .A3(new_n260), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT25), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n221), .A2(new_n271), .ZN(new_n437));
  INV_X1    g0237(.A(G257), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G1698), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n328), .A2(new_n437), .A3(new_n330), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G294), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT80), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT80), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G294), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n444), .A3(G33), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT81), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT81), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n274), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G41), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n212), .B(G45), .C1(new_n451), .C2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT74), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G1), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT74), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n457), .B2(G41), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n451), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n460), .A2(G274), .A3(new_n280), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n452), .A2(KEYINPUT74), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n456), .B1(new_n455), .B2(new_n458), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G264), .A3(new_n280), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n450), .A2(G179), .A3(new_n465), .A4(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n475), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n436), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n471), .A2(new_n475), .A3(new_n472), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n471), .B2(new_n472), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n436), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n331), .B1(G264), .B2(G1698), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n438), .B2(G1698), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n274), .C1(G303), .C2(new_n269), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n274), .B1(new_n460), .B2(new_n464), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(G270), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n488), .B2(G270), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n487), .B(new_n465), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n263), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(G20), .B1(G33), .B2(G283), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(G33), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n258), .B(new_n497), .C1(new_n213), .C2(G116), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT20), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  OAI221_X1 g0301(.A(new_n494), .B1(new_n493), .B2(new_n431), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n492), .A2(new_n502), .A3(G169), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT21), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n492), .A2(G200), .ZN(new_n506));
  INV_X1    g0306(.A(new_n502), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(new_n284), .C2(new_n492), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n492), .A2(new_n301), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n502), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n492), .A2(new_n502), .A3(KEYINPUT21), .A4(G169), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n505), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n429), .A2(new_n433), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n450), .A2(new_n469), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(G190), .A3(new_n465), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n470), .A2(G200), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n435), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g0318(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n328), .A2(new_n330), .A3(new_n271), .ZN(new_n520));
  OAI21_X1  g0320(.A(G244), .B1(KEYINPUT73), .B2(KEYINPUT4), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n221), .A2(new_n271), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n269), .A2(new_n523), .B1(G33), .B2(G283), .ZN(new_n524));
  INV_X1    g0324(.A(new_n521), .ZN(new_n525));
  INV_X1    g0325(.A(new_n519), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n269), .A2(new_n271), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n274), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n468), .A2(G257), .A3(new_n280), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(new_n301), .A3(new_n465), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  AND2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n417), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n213), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n359), .A2(new_n360), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G107), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n254), .A2(new_n218), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n257), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n262), .A2(G97), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n432), .B2(G97), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n531), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AOI221_X4 g0346(.A(new_n277), .B1(new_n462), .B2(new_n463), .C1(new_n453), .C2(new_n459), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n280), .A2(new_n547), .B1(new_n488), .B2(G257), .ZN(new_n548));
  AOI21_X1  g0348(.A(G169), .B1(new_n548), .B2(new_n529), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n518), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n529), .A2(new_n465), .A3(new_n530), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n290), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n540), .B(new_n537), .C1(new_n538), .C2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n544), .B1(new_n553), .B2(new_n257), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT76), .A4(new_n531), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n554), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(G200), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n284), .C2(new_n551), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n226), .A2(new_n271), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n219), .A2(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n328), .A2(new_n560), .A3(new_n330), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G116), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n566), .A2(new_n567), .A3(new_n280), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n221), .B1(new_n454), .B2(G1), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n455), .A2(new_n277), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n280), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n290), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n303), .A2(new_n262), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n213), .B1(new_n325), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n220), .A2(new_n496), .A3(new_n417), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n269), .A2(new_n213), .A3(G68), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(KEYINPUT78), .A3(new_n577), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n575), .B1(new_n314), .B2(new_n496), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n574), .B1(new_n584), .B2(new_n258), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n432), .A2(new_n303), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n567), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n274), .A3(new_n565), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n301), .A3(new_n571), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n573), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n568), .B2(new_n572), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n431), .A2(new_n220), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n574), .B(new_n593), .C1(new_n584), .C2(new_n258), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n589), .A2(G190), .A3(new_n571), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n556), .A2(new_n559), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n484), .A2(new_n512), .A3(new_n517), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n416), .A2(new_n600), .ZN(G372));
  INV_X1    g0401(.A(new_n292), .ZN(new_n602));
  INV_X1    g0402(.A(new_n310), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n344), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n342), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n396), .A3(new_n400), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n408), .A2(KEYINPUT85), .A3(new_n401), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT85), .B1(new_n408), .B2(new_n401), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT18), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n410), .A3(new_n607), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n602), .B1(new_n614), .B2(new_n288), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n550), .A2(new_n555), .A3(new_n591), .A4(new_n596), .ZN(new_n616));
  XNOR2_X1  g0416(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n552), .A2(new_n554), .A3(new_n531), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n597), .A2(new_n618), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n616), .A2(new_n617), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n517), .A2(new_n556), .A3(new_n559), .A4(new_n598), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n436), .A2(new_n473), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n505), .A2(new_n622), .A3(new_n510), .A4(new_n511), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n591), .B(new_n620), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n415), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n615), .A2(new_n625), .ZN(G369));
  AND2_X1   g0426(.A1(new_n484), .A2(new_n517), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n260), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n261), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT86), .Z(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n436), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT87), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n636), .A2(KEYINPUT87), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n627), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n481), .A2(new_n436), .A3(new_n635), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n502), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n512), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n505), .A2(new_n510), .A3(new_n511), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(new_n635), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n627), .A2(new_n637), .A3(new_n638), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n635), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n436), .A2(new_n473), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n648), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n214), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G1), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n577), .A2(G116), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(new_n210), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT29), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n482), .B1(new_n481), .B2(new_n436), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n482), .A2(new_n436), .A3(new_n474), .A4(new_n476), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n645), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n517), .A2(new_n556), .A3(new_n559), .A4(new_n598), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n616), .A2(new_n617), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n619), .A2(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n591), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n616), .A2(new_n617), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n673));
  INV_X1    g0473(.A(new_n591), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT89), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n667), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n662), .B1(new_n676), .B2(new_n651), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n624), .A2(new_n651), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(KEYINPUT29), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n488), .A2(G270), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT79), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n488), .A2(new_n489), .A3(G270), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n683), .A2(new_n684), .B1(new_n280), .B2(new_n547), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(G179), .A3(new_n487), .A4(new_n514), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n589), .A2(new_n571), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n551), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n681), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n514), .A4(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n551), .A2(new_n470), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n492), .A2(new_n301), .A3(new_n687), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT88), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n492), .A2(new_n696), .A3(new_n301), .A4(new_n687), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n693), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n635), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT31), .B(new_n635), .C1(new_n692), .C2(new_n698), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n701), .B(new_n702), .C1(new_n600), .C2(new_n635), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n680), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n661), .B1(new_n706), .B2(G1), .ZN(G364));
  AOI21_X1  g0507(.A(new_n206), .B1(G20), .B2(new_n290), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G179), .A2(G200), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT93), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n213), .A2(G190), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  XOR2_X1   g0514(.A(KEYINPUT94), .B(G159), .Z(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT32), .ZN(new_n717));
  INV_X1    g0517(.A(G200), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G179), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT95), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(G20), .A3(G190), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G87), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n712), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n723), .B(new_n269), .C1(new_n417), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(G20), .A2(G179), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n728), .A2(new_n284), .A3(G200), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n225), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n717), .A2(new_n725), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n284), .A3(new_n718), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(KEYINPUT91), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(KEYINPUT91), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n728), .A2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n718), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n738), .A2(G77), .B1(G50), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n728), .A2(G190), .A3(new_n718), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n362), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n732), .B1(new_n733), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n711), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n744), .B1(new_n733), .B2(new_n743), .C1(new_n496), .C2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n730), .A2(new_n749), .B1(new_n750), .B2(new_n742), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT96), .B(G326), .Z(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(new_n740), .B1(new_n714), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n724), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n442), .A2(new_n444), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n751), .B(new_n755), .C1(new_n757), .C2(new_n746), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n269), .B1(new_n722), .B2(G303), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n738), .A2(G311), .B1(new_n759), .B2(KEYINPUT97), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n758), .B(new_n760), .C1(KEYINPUT97), .C2(new_n759), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n709), .B1(new_n748), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n708), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n655), .A2(new_n269), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n210), .A2(G45), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n243), .C2(new_n454), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n655), .A2(new_n331), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G355), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n769), .B(new_n771), .C1(G116), .C2(new_n214), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n762), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n765), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n646), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n658), .B1(G45), .B2(new_n628), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n646), .A2(G330), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n647), .A2(new_n777), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n775), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(G396));
  NOR2_X1   g0580(.A1(new_n310), .A2(new_n635), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n635), .A2(new_n309), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n350), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n310), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n678), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n781), .B1(new_n310), .B2(new_n784), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n624), .A2(new_n651), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(new_n704), .Z(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n777), .ZN(new_n792));
  INV_X1    g0592(.A(new_n742), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G137), .A2(new_n740), .B1(new_n793), .B2(G143), .ZN(new_n794));
  INV_X1    g0594(.A(new_n715), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n252), .B2(new_n730), .C1(new_n737), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT34), .ZN(new_n797));
  INV_X1    g0597(.A(new_n724), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G68), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n269), .B1(new_n713), .B2(new_n800), .C1(new_n721), .C2(new_n202), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G58), .B2(new_n746), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n797), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n740), .ZN(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n747), .A2(new_n496), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n331), .B1(new_n724), .B2(new_n220), .C1(new_n417), .C2(new_n721), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n713), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n730), .A2(new_n754), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n806), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n493), .B2(new_n737), .C1(new_n441), .C2(new_n742), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n709), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n708), .A2(new_n763), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G77), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n776), .C1(new_n764), .C2(new_n788), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n792), .A2(new_n818), .ZN(G384));
  NOR3_X1   g0619(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n820));
  OAI211_X1 g0620(.A(KEYINPUT100), .B(new_n344), .C1(new_n820), .C2(new_n322), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n821), .A2(new_n323), .A3(new_n635), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n635), .A2(new_n323), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n342), .A2(KEYINPUT100), .A3(new_n344), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n786), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n633), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n372), .A2(new_n258), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT16), .B1(new_n370), .B2(new_n371), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n386), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n414), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n405), .A2(new_n408), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n405), .A2(new_n826), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT37), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n392), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n412), .A2(new_n633), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n397), .B1(new_n835), .B2(new_n829), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n830), .A2(KEYINPUT38), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n830), .B2(new_n837), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n703), .B(new_n825), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT40), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n825), .A2(KEYINPUT40), .A3(new_n703), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(KEYINPUT103), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n392), .B(KEYINPUT102), .Z(new_n846));
  NAND4_X1  g0646(.A1(new_n846), .A2(new_n611), .A3(new_n607), .A4(new_n832), .ZN(new_n847));
  AOI211_X1 g0647(.A(KEYINPUT37), .B(new_n397), .C1(new_n405), .C2(new_n408), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(KEYINPUT37), .B1(new_n832), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n394), .A2(new_n395), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n832), .B1(new_n613), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n845), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT103), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n830), .A2(new_n853), .A3(KEYINPUT38), .A4(new_n837), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n844), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n841), .A2(new_n842), .B1(new_n843), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT104), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n415), .A2(new_n703), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(G330), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n830), .A2(new_n837), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n845), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(KEYINPUT39), .A3(new_n838), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n342), .A2(new_n635), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n789), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n822), .A2(new_n824), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(new_n839), .C2(new_n840), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT101), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n610), .A2(new_n612), .A3(new_n633), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n415), .B1(new_n677), .B2(new_n679), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n615), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n877), .B(new_n879), .Z(new_n880));
  XNOR2_X1  g0680(.A(new_n860), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n212), .B2(new_n628), .ZN(new_n882));
  INV_X1    g0682(.A(new_n209), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n535), .A2(new_n536), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n493), .B1(new_n884), .B2(KEYINPUT35), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n883), .B(new_n885), .C1(KEYINPUT35), .C2(new_n884), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT36), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n363), .A2(new_n210), .A3(new_n218), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT98), .Z(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(G50), .B2(new_n225), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(G1), .A3(new_n260), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n882), .A2(new_n887), .A3(new_n891), .ZN(G367));
  OAI211_X1 g0692(.A(new_n556), .B(new_n559), .C1(new_n557), .C2(new_n651), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n651), .A2(new_n618), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n648), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n651), .A2(new_n594), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n674), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n597), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT106), .Z(new_n902));
  XNOR2_X1  g0702(.A(new_n897), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n650), .A2(new_n893), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT42), .Z(new_n906));
  NAND3_X1  g0706(.A1(new_n896), .A2(new_n478), .A3(new_n483), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n635), .B1(new_n907), .B2(new_n556), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n903), .B(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n656), .B(KEYINPUT41), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n895), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT107), .B1(new_n653), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n650), .A2(new_n915), .A3(new_n652), .A4(new_n895), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT45), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n653), .A2(new_n913), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT44), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(KEYINPUT45), .A3(new_n916), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(KEYINPUT44), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n919), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n648), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  INV_X1    g0726(.A(new_n648), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(new_n921), .A4(new_n919), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n641), .A2(new_n649), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n650), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(new_n647), .Z(new_n931));
  NAND4_X1  g0731(.A1(new_n925), .A2(new_n928), .A3(new_n931), .A4(new_n706), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n912), .B1(new_n932), .B2(new_n706), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n212), .B1(new_n628), .B2(G45), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n910), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT46), .B1(new_n722), .B2(G116), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G303), .B2(new_n793), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n417), .B2(new_n747), .C1(new_n808), .C2(new_n804), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n722), .A2(KEYINPUT46), .A3(G116), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n714), .A2(G317), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n729), .A2(new_n757), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n940), .A2(new_n331), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n737), .A2(new_n754), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n724), .A2(new_n496), .ZN(new_n945));
  NOR4_X1   g0745(.A1(new_n939), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n729), .A2(new_n715), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n746), .A2(G68), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n740), .A2(G143), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n252), .C2(new_n742), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n331), .B1(new_n722), .B2(G58), .ZN(new_n951));
  INV_X1    g0751(.A(G137), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n951), .B1(new_n218), .B2(new_n724), .C1(new_n952), .C2(new_n713), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n950), .B(new_n953), .C1(G50), .C2(new_n738), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n946), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  AOI21_X1  g0756(.A(new_n777), .B1(new_n956), .B2(new_n708), .ZN(new_n957));
  INV_X1    g0757(.A(new_n303), .ZN(new_n958));
  INV_X1    g0758(.A(new_n767), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n766), .B1(new_n214), .B2(new_n958), .C1(new_n239), .C2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(new_n774), .C2(new_n900), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n936), .A2(new_n961), .ZN(G387));
  OR2_X1    g0762(.A1(new_n931), .A2(new_n706), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n931), .A2(new_n706), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n656), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n959), .B1(new_n236), .B2(G45), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n659), .B2(new_n770), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n248), .A2(new_n202), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n659), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n969), .B(new_n454), .C1(KEYINPUT50), .C2(new_n968), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G68), .B2(G77), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n967), .A2(new_n971), .B1(G107), .B2(new_n214), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n777), .B1(new_n972), .B2(new_n766), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n331), .B1(new_n724), .B2(new_n493), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT108), .B(G322), .Z(new_n975));
  AOI22_X1  g0775(.A1(new_n740), .A2(new_n975), .B1(new_n729), .B2(G311), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n976), .B1(new_n977), .B2(new_n742), .C1(new_n737), .C2(new_n805), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n754), .B2(new_n747), .C1(new_n756), .C2(new_n721), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT49), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n974), .B(new_n982), .C1(new_n752), .C2(new_n714), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n747), .A2(new_n958), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n248), .B2(new_n729), .ZN(new_n985));
  INV_X1    g0785(.A(G159), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n986), .B2(new_n804), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n737), .A2(new_n225), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n945), .A2(new_n331), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n722), .A2(G77), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n252), .C2(new_n713), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n742), .A2(new_n202), .ZN(new_n992));
  NOR4_X1   g0792(.A1(new_n987), .A2(new_n988), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n983), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT109), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n973), .B1(new_n641), .B2(new_n774), .C1(new_n996), .C2(new_n709), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n931), .A2(new_n935), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n965), .A2(new_n997), .A3(new_n998), .ZN(G393));
  NAND2_X1  g0799(.A1(new_n925), .A2(new_n928), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n964), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(new_n656), .A3(new_n932), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n925), .A2(new_n928), .A3(new_n935), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n896), .A2(new_n774), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT110), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n766), .B1(new_n496), .B2(new_n214), .C1(new_n246), .C2(new_n959), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(KEYINPUT110), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n747), .A2(new_n218), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n269), .B1(new_n724), .B2(new_n220), .C1(new_n225), .C2(new_n721), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G50), .C2(new_n729), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n714), .A2(G143), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n804), .A2(new_n252), .B1(new_n986), .B2(new_n742), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT51), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n248), .A2(new_n738), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1010), .A2(new_n1011), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n804), .A2(new_n977), .B1(new_n808), .B2(new_n742), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n746), .A2(G116), .B1(new_n729), .B2(G303), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT111), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n331), .B1(new_n724), .B2(new_n417), .C1(new_n754), .C2(new_n721), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n738), .B2(G294), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n714), .A2(new_n975), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1016), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n777), .B1(new_n1025), .B2(new_n708), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1002), .A2(new_n1003), .A3(new_n1027), .ZN(G390));
  NAND3_X1  g0828(.A1(new_n415), .A2(G330), .A3(new_n703), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n878), .A2(new_n615), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n825), .A2(G330), .A3(new_n703), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n703), .A2(G330), .A3(new_n788), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n871), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n676), .A2(new_n651), .A3(new_n785), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n782), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1031), .B(new_n1034), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(new_n1031), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n870), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1030), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1035), .A2(new_n782), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT112), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n871), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n866), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n855), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n862), .A2(new_n865), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n870), .A2(new_n871), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n1047), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1031), .A2(KEYINPUT113), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1050), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1041), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1055), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1048), .B1(new_n1060), .B2(new_n871), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n862), .A2(new_n865), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1050), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1030), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1058), .A2(new_n656), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n723), .A2(new_n331), .A3(new_n799), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1008), .B1(G283), .B2(new_n740), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n493), .B2(new_n742), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G294), .C2(new_n714), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n496), .B2(new_n737), .C1(new_n417), .C2(new_n730), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT115), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n747), .A2(new_n986), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n804), .A2(new_n1078), .B1(new_n800), .B2(new_n742), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(G137), .C2(new_n729), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n722), .A2(G150), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT53), .Z(new_n1082));
  AOI21_X1  g0882(.A(new_n331), .B1(new_n714), .B2(G125), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1084), .B1(new_n202), .B2(new_n724), .C1(new_n737), .C2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT114), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n708), .B1(new_n1076), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n776), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1051), .B2(new_n763), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n248), .B2(new_n815), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1070), .A2(new_n935), .B1(KEYINPUT116), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(KEYINPUT116), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1069), .A2(new_n1093), .A3(new_n1094), .ZN(G378));
  NAND2_X1  g0895(.A1(new_n841), .A2(new_n842), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n843), .A2(new_n855), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(G330), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n288), .A2(new_n292), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT55), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n826), .A2(new_n266), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT56), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1100), .B(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n856), .B2(G330), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n877), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n872), .A2(new_n874), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT101), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n856), .A2(G330), .A3(new_n1103), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n867), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n934), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1104), .A2(new_n763), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n814), .A2(new_n202), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n798), .A2(G58), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n990), .A2(new_n1118), .A3(new_n451), .A4(new_n331), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n948), .B1(new_n417), .B2(new_n742), .C1(new_n496), .C2(new_n730), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(G283), .C2(new_n714), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n493), .B2(new_n804), .C1(new_n958), .C2(new_n737), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT58), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(G33), .A2(G41), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT117), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1125), .B(new_n202), .C1(G41), .C2(new_n269), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n746), .A2(G150), .B1(new_n740), .B2(G125), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT118), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n730), .A2(new_n800), .B1(new_n721), .B2(new_n1086), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n738), .B2(G137), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(new_n1078), .C2(new_n742), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n798), .A2(new_n715), .B1(new_n714), .B2(G124), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1123), .B(new_n1126), .C1(new_n1125), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n777), .B1(new_n1136), .B2(new_n708), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1116), .A2(new_n1117), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1115), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1107), .A2(new_n1114), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1067), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1142));
  OAI211_X1 g0942(.A(KEYINPUT57), .B(new_n1141), .C1(new_n1142), .C2(new_n1030), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n656), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1058), .A2(new_n1066), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT57), .B1(new_n1145), .B2(new_n1141), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1140), .B1(new_n1144), .B2(new_n1146), .ZN(G375));
  NOR2_X1   g0947(.A1(new_n871), .A2(new_n764), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n331), .B1(new_n713), .B2(new_n805), .C1(new_n724), .C2(new_n218), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n984), .B1(G116), .B2(new_n729), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n754), .B2(new_n742), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(G97), .C2(new_n722), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n417), .B2(new_n737), .C1(new_n441), .C2(new_n804), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1118), .B(new_n269), .C1(new_n986), .C2(new_n721), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n747), .A2(new_n202), .B1(new_n952), .B2(new_n742), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n713), .A2(new_n1078), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n730), .A2(new_n1086), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n800), .B2(new_n804), .C1(new_n252), .C2(new_n737), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n709), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n815), .A2(G68), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1148), .A2(new_n777), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1065), .B2(new_n935), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1038), .A2(new_n1040), .A3(new_n1030), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n911), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1165), .B2(new_n1041), .ZN(G381));
  OAI21_X1  g0966(.A(new_n1141), .B1(new_n1142), .B2(new_n1030), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n656), .A3(new_n1143), .ZN(new_n1170));
  INV_X1    g0970(.A(G378), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1140), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1172), .A2(G384), .A3(G381), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(G387), .A2(G390), .A3(G396), .A4(G393), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(G407));
  OAI211_X1 g0975(.A(G407), .B(G213), .C1(G343), .C2(new_n1172), .ZN(G409));
  INV_X1    g0976(.A(G390), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(G387), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(G390), .A2(new_n936), .A3(new_n961), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(KEYINPUT121), .A3(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(G393), .B(G396), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT121), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(G387), .A2(new_n1177), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1178), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(G387), .A2(new_n1177), .A3(KEYINPUT122), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1179), .B(KEYINPUT123), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1185), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1141), .A2(new_n935), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(KEYINPUT119), .A3(new_n1138), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT119), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1115), .B2(new_n1139), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1058), .A2(new_n1066), .B1(new_n1114), .B2(new_n1107), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1193), .A2(new_n1195), .B1(new_n1196), .B2(new_n911), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1197), .A2(new_n1171), .B1(G213), .B2(new_n634), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(G375), .A2(G378), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT60), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1067), .B(new_n656), .C1(new_n1200), .C2(new_n1164), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1164), .A2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1163), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G384), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT120), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT120), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(new_n1208), .A3(new_n1204), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1198), .A2(new_n1199), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT63), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(KEYINPUT63), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1191), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT61), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n634), .A2(G213), .A3(G2897), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1210), .B(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1216), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1215), .B(new_n1222), .C1(KEYINPUT124), .C2(new_n1191), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT124), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT62), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1212), .A2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT125), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1198), .A2(new_n1199), .A3(new_n1211), .A4(KEYINPUT62), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(KEYINPUT125), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1225), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1223), .B1(new_n1231), .B2(new_n1191), .ZN(G405));
  NOR2_X1   g1032(.A1(G375), .A2(G378), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1171), .B1(new_n1170), .B2(new_n1140), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT126), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT127), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1211), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1199), .B2(new_n1172), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT127), .B1(new_n1239), .B2(new_n1210), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1233), .A2(new_n1234), .A3(KEYINPUT126), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1237), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1191), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1191), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1236), .B1(new_n1235), .B2(new_n1211), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n1210), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1237), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1246), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1245), .A2(new_n1251), .ZN(G402));
endmodule


