//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n475), .A2(KEYINPUT66), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n465), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n474), .B2(new_n477), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n468), .B2(new_n469), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n463), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n475), .B2(new_n476), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n465), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT67), .B1(new_n503), .B2(KEYINPUT68), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT5), .B1(new_n503), .B2(KEYINPUT67), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(KEYINPUT67), .B(KEYINPUT5), .C1(new_n503), .C2(KEYINPUT68), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n506), .A2(G88), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n506), .A2(G62), .A3(new_n507), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G166));
  AND2_X1   g092(.A1(new_n506), .A2(new_n507), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT70), .B(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n508), .A2(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT69), .B(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n523), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(new_n522), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n506), .A2(new_n507), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n520), .A2(G90), .B1(G52), .B2(new_n523), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n532), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n520), .A2(G81), .B1(G43), .B2(new_n523), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G860), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n520), .A2(G91), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n523), .A2(G53), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n553), .B(KEYINPUT9), .C1(new_n511), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT73), .B(G65), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n506), .A2(new_n507), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n559), .B1(new_n563), .B2(G651), .ZN(new_n564));
  AOI211_X1 g139(.A(KEYINPUT74), .B(new_n513), .C1(new_n561), .C2(new_n562), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n552), .B(new_n558), .C1(new_n564), .C2(new_n565), .ZN(G299));
  NAND2_X1  g141(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n535), .A2(new_n536), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G301));
  INV_X1    g146(.A(new_n512), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n514), .A2(new_n515), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G303));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n513), .B1(new_n532), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(G49), .B2(new_n523), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n520), .A2(G87), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(new_n520), .B2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n523), .A2(G48), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n506), .A2(G86), .A3(new_n507), .A4(new_n508), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n506), .A2(G61), .A3(new_n507), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT77), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n513), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n520), .A2(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n511), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n518), .A2(G60), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n513), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(KEYINPUT78), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n532), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT79), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n608), .B(new_n604), .C1(new_n532), .C2(new_n605), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(G651), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n506), .A2(G92), .A3(new_n507), .A4(new_n508), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n611), .A2(new_n614), .B1(G54), .B2(new_n523), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n602), .B1(new_n603), .B2(new_n617), .ZN(G284));
  AOI21_X1  g193(.A(new_n602), .B1(new_n603), .B2(new_n617), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n558), .A2(new_n552), .ZN(new_n621));
  INV_X1    g196(.A(new_n564), .ZN(new_n622));
  INV_X1    g197(.A(new_n565), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(new_n624), .B2(G868), .ZN(G280));
  XNOR2_X1  g200(.A(G280), .B(KEYINPUT80), .ZN(G297));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n616), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(new_n544), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT81), .B1(new_n629), .B2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n616), .A2(new_n627), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  MUX2_X1   g207(.A(KEYINPUT81), .B(new_n630), .S(new_n632), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n479), .A2(G135), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(G111), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(G2105), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n482), .B2(G123), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2096), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  NOR2_X1   g244(.A1(G2072), .A2(G2078), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(KEYINPUT85), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(KEYINPUT85), .ZN(new_n674));
  INV_X1    g249(.A(new_n669), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n671), .B(KEYINPUT17), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  INV_X1    g254(.A(new_n667), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n669), .A2(new_n680), .A3(new_n671), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n669), .A2(new_n667), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n679), .B(new_n682), .C1(new_n676), .C2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n691), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT20), .Z(new_n695));
  AOI211_X1 g270(.A(new_n693), .B(new_n695), .C1(new_n688), .C2(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT88), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT87), .Z(new_n699));
  XOR2_X1   g274(.A(G1981), .B(G1986), .Z(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n697), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G19), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n629), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1341), .ZN(new_n708));
  INV_X1    g283(.A(G2067), .ZN(new_n709));
  INV_X1    g284(.A(G104), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n710), .A2(new_n465), .A3(KEYINPUT92), .ZN(new_n711));
  AOI21_X1  g286(.A(KEYINPUT92), .B1(new_n710), .B2(new_n465), .ZN(new_n712));
  OAI221_X1 g287(.A(G2104), .B1(G116), .B2(new_n465), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G140), .ZN(new_n714));
  INV_X1    g289(.A(G128), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n713), .B1(new_n478), .B2(new_n714), .C1(new_n715), .C2(new_n481), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G26), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT93), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n709), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n717), .A2(new_n709), .A3(new_n721), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n708), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n616), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G4), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n724), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n718), .A2(G35), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G162), .B2(new_n718), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G2090), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G33), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT95), .Z(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n465), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G139), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT25), .Z(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT97), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G2072), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n736), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n748), .A2(G2072), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n735), .A2(G2090), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n730), .A2(new_n731), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n705), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n705), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G1961), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n718), .A2(G32), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT102), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G141), .B2(new_n479), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT101), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n482), .B2(G129), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n758), .B1(new_n767), .B2(new_n718), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n757), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n718), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n718), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G2078), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G2078), .ZN(new_n776));
  INV_X1    g351(.A(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(KEYINPUT30), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n775), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G1961), .B2(new_n756), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n642), .A2(G29), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n718), .B1(new_n786), .B2(G34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(G34), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT99), .Z(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G29), .B2(G160), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT100), .B(G2084), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n705), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n705), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n784), .A2(new_n785), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n705), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n624), .B2(new_n705), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1956), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n772), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n732), .A2(new_n753), .A3(new_n754), .A4(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G23), .B(G288), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n705), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n705), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1971), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n705), .A2(G6), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n591), .B2(new_n705), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT32), .B(G1981), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT90), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n809), .A2(new_n814), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n479), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n482), .A2(G119), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n465), .A2(G107), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G25), .B(new_n828), .S(G29), .Z(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n705), .A2(G24), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n599), .B2(new_n705), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT89), .B(G1986), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n822), .A2(new_n823), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n822), .A2(new_n840), .A3(new_n823), .A4(new_n837), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n806), .B1(new_n839), .B2(new_n841), .ZN(G311));
  XNOR2_X1  g417(.A(G311), .B(KEYINPUT103), .ZN(G150));
  NAND2_X1  g418(.A1(new_n610), .A2(new_n615), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n627), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n532), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G651), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n523), .A2(G55), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n506), .A2(G93), .A3(new_n507), .A4(new_n508), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n544), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n857), .A2(new_n542), .A3(new_n851), .A4(new_n543), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n847), .B(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n545), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n852), .A2(new_n855), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n545), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(G145));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n496), .B2(new_n499), .ZN(new_n869));
  OAI211_X1 g444(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n469), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(KEYINPUT106), .C1(new_n497), .C2(new_n498), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n494), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n716), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n716), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n767), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n747), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n747), .A2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n875), .A2(new_n766), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n879), .B(new_n747), .C1(new_n877), .C2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n479), .A2(G142), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n482), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n465), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n647), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(new_n828), .Z(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n884), .A2(new_n885), .A3(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G160), .B(KEYINPUT105), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n486), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n643), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n900), .A3(new_n896), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n907));
  NAND2_X1  g482(.A1(G303), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(G166), .A2(KEYINPUT109), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n908), .A2(G305), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G305), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G288), .B(new_n599), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  NOR2_X1   g491(.A1(G290), .A2(G288), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n579), .B(new_n580), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n599), .B1(new_n918), .B2(new_n578), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n913), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(KEYINPUT110), .A3(new_n914), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n856), .A2(new_n858), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n631), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n624), .A2(new_n844), .ZN(new_n927));
  NAND3_X1  g502(.A1(G299), .A2(new_n610), .A3(new_n615), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT41), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n624), .A2(new_n844), .A3(KEYINPUT108), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n928), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n930), .B1(new_n937), .B2(new_n926), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n924), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G868), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g516(.A(new_n940), .B1(G868), .B2(new_n864), .ZN(G331));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  AOI21_X1  g518(.A(G286), .B1(new_n567), .B2(new_n569), .ZN(new_n944));
  NOR2_X1   g519(.A1(G171), .A2(G168), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n925), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT112), .B(new_n925), .C1(new_n944), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n570), .A2(G168), .ZN(new_n951));
  INV_X1    g526(.A(new_n945), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n859), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n929), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n931), .ZN(new_n956));
  INV_X1    g531(.A(new_n934), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT108), .B1(new_n624), .B2(new_n844), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n624), .A2(new_n844), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n960), .B2(KEYINPUT41), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n953), .A2(new_n946), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n953), .A2(new_n946), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT111), .B1(new_n937), .B2(new_n965), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n923), .B(new_n955), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n953), .A2(new_n929), .A3(new_n946), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n948), .A2(new_n953), .A3(new_n949), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n933), .A2(KEYINPUT41), .A3(new_n928), .A4(new_n934), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n929), .A2(new_n936), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n923), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n903), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n955), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n962), .B1(new_n961), .B2(new_n963), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n937), .A2(new_n965), .A3(KEYINPUT111), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n975), .B(new_n978), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n970), .A2(new_n973), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n968), .ZN(new_n983));
  AOI21_X1  g558(.A(G37), .B1(new_n983), .B2(new_n923), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n977), .A2(KEYINPUT43), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n955), .B1(new_n964), .B2(new_n966), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n903), .B1(new_n990), .B2(new_n975), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n943), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n991), .B2(new_n967), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n981), .A2(new_n984), .A3(new_n988), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n994), .A2(new_n943), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(G397));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n872), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n872), .A2(KEYINPUT117), .A3(new_n1000), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G160), .A2(G40), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n501), .A2(new_n1000), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(KEYINPUT50), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2084), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT122), .B1(new_n1012), .B2(new_n1007), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n872), .A2(KEYINPUT117), .A3(new_n1000), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT117), .B1(new_n872), .B2(new_n1000), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1007), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1013), .A2(new_n1014), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1011), .B1(new_n1022), .B2(new_n798), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n999), .B1(new_n1023), .B2(G168), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1014), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n798), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1011), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G286), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n998), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT51), .B(new_n999), .C1(new_n1023), .C2(G168), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT62), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1027), .A2(G168), .A3(new_n1028), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1023), .A2(G168), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT51), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1024), .A2(new_n998), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1016), .A2(new_n1017), .A3(new_n1007), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n999), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n918), .A2(G1976), .A3(new_n578), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  INV_X1    g623(.A(new_n586), .ZN(new_n1049));
  INV_X1    g624(.A(new_n590), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n586), .A2(new_n590), .A3(G1981), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT118), .B(new_n1047), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT118), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1042), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1020), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1043), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1046), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n512), .B2(new_n516), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT55), .ZN(new_n1062));
  INV_X1    g637(.A(G2090), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1006), .A2(new_n1009), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1020), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT116), .B(G1971), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n999), .B(new_n1062), .C1(new_n1064), .C2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1060), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1062), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1004), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1007), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT50), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT120), .A3(new_n1020), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT121), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1075), .A2(new_n1063), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n999), .B1(new_n1080), .B2(new_n1069), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1071), .B1(new_n1072), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G2078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1013), .A2(new_n1014), .A3(new_n1021), .A4(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1067), .A2(G2078), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1010), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n570), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1082), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1033), .A2(new_n1040), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT119), .Z(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1042), .B1(new_n1096), .B2(new_n1052), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1070), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1060), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1029), .A2(G8), .A3(G168), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1100), .B1(new_n1082), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1100), .B1(new_n1104), .B2(new_n1062), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1071), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1099), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1020), .A2(new_n1066), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1065), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1075), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(KEYINPUT123), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT57), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1348), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1057), .A2(G2067), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n616), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1124));
  AND4_X1   g699(.A1(KEYINPUT61), .A2(new_n1124), .A3(new_n1117), .A4(new_n1111), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT125), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n616), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n616), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n844), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(KEYINPUT60), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  INV_X1    g711(.A(G1996), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1020), .A2(new_n1065), .A3(new_n1137), .A4(new_n1066), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT58), .B(G1341), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1041), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT124), .B(new_n1138), .C1(new_n1041), .C2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1136), .B1(new_n1144), .B2(new_n629), .ZN(new_n1145));
  AOI211_X1 g720(.A(KEYINPUT59), .B(new_n544), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1132), .B(new_n1135), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1129), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1115), .A2(new_n1149), .A3(new_n1117), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1126), .B1(new_n1150), .B2(new_n1119), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1123), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT45), .B1(new_n872), .B2(new_n1000), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1153), .A2(new_n1083), .A3(G2078), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1086), .A2(new_n1083), .B1(new_n1109), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(G301), .A3(new_n1089), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT54), .B1(new_n1091), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n1082), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT126), .B1(new_n1090), .B2(new_n570), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1160), .A2(new_n1161), .A3(G301), .A4(new_n1085), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1155), .A2(new_n1089), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(G171), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1158), .B(new_n1167), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1093), .B(new_n1108), .C1(new_n1152), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1020), .A2(new_n1153), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n716), .B(G2067), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT115), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n766), .A2(G1996), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1171), .A2(G1996), .A3(new_n766), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT114), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n828), .B(new_n830), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1175), .B(new_n1177), .C1(new_n1170), .C2(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  NAND2_X1  g755(.A1(G290), .A2(G1986), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1170), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1169), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1180), .A2(new_n1170), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT127), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT48), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT47), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1171), .B1(new_n1173), .B2(new_n766), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1171), .A2(new_n1137), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT46), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1188), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n1187), .A2(new_n1179), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n828), .A2(new_n831), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1175), .A2(new_n1196), .A3(new_n1177), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n716), .A2(G2067), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1170), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1184), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g776(.A1(new_n994), .A2(new_n995), .ZN(new_n1203));
  NOR4_X1   g777(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n1203), .A2(new_n905), .A3(new_n1204), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


