

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736;

  XNOR2_X1 U363 ( .A(n527), .B(n526), .ZN(n588) );
  NAND2_X1 U364 ( .A1(n525), .A2(n524), .ZN(n527) );
  BUF_X1 U365 ( .A(n516), .Z(n341) );
  XNOR2_X1 U366 ( .A(n342), .B(n519), .ZN(n674) );
  NAND2_X1 U367 ( .A1(n393), .A2(n350), .ZN(n342) );
  OR2_X1 U368 ( .A1(n620), .A2(G902), .ZN(n400) );
  XNOR2_X1 U369 ( .A(n714), .B(n418), .ZN(n504) );
  XNOR2_X1 U370 ( .A(n413), .B(n411), .ZN(n714) );
  AND2_X1 U371 ( .A1(n736), .A2(n632), .ZN(n587) );
  XNOR2_X1 U372 ( .A(G116), .B(KEYINPUT73), .ZN(n376) );
  XNOR2_X1 U373 ( .A(G119), .B(G110), .ZN(n458) );
  XNOR2_X1 U374 ( .A(n392), .B(G131), .ZN(n488) );
  XNOR2_X2 U375 ( .A(n473), .B(n472), .ZN(n649) );
  XNOR2_X2 U376 ( .A(n608), .B(n354), .ZN(n372) );
  NOR2_X2 U377 ( .A1(n569), .A2(n571), .ZN(n500) );
  XNOR2_X2 U378 ( .A(KEYINPUT10), .B(n461), .ZN(n727) );
  XNOR2_X2 U379 ( .A(G146), .B(KEYINPUT68), .ZN(n392) );
  XNOR2_X1 U380 ( .A(n594), .B(n593), .ZN(n629) );
  NAND2_X1 U381 ( .A1(n387), .A2(n386), .ZN(n596) );
  INV_X2 U382 ( .A(G953), .ZN(n391) );
  XNOR2_X1 U383 ( .A(KEYINPUT84), .B(G143), .ZN(n422) );
  XNOR2_X1 U384 ( .A(n497), .B(KEYINPUT107), .ZN(n499) );
  AND2_X1 U385 ( .A1(n386), .A2(n389), .ZN(n385) );
  AND2_X1 U386 ( .A1(n388), .A2(n347), .ZN(n387) );
  OR2_X2 U387 ( .A1(n545), .A2(n346), .ZN(n386) );
  NOR2_X1 U388 ( .A1(n667), .A2(n668), .ZN(n410) );
  XNOR2_X1 U389 ( .A(n494), .B(KEYINPUT99), .ZN(n556) );
  XNOR2_X1 U390 ( .A(n356), .B(G478), .ZN(n528) );
  XOR2_X1 U391 ( .A(n701), .B(KEYINPUT59), .Z(n702) );
  XNOR2_X1 U392 ( .A(n401), .B(n726), .ZN(n620) );
  XNOR2_X1 U393 ( .A(n405), .B(n404), .ZN(n701) );
  XNOR2_X1 U394 ( .A(n504), .B(n503), .ZN(n401) );
  XNOR2_X1 U395 ( .A(n490), .B(n406), .ZN(n405) );
  XNOR2_X1 U396 ( .A(n422), .B(n421), .ZN(n440) );
  INV_X1 U397 ( .A(G140), .ZN(n501) );
  XNOR2_X1 U398 ( .A(G107), .B(G110), .ZN(n414) );
  XNOR2_X1 U399 ( .A(KEYINPUT3), .B(G113), .ZN(n375) );
  AND2_X1 U400 ( .A1(n372), .A2(n609), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n417), .B(n414), .ZN(n413) );
  BUF_X1 U402 ( .A(n664), .Z(n344) );
  INV_X1 U403 ( .A(n571), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n410), .B(KEYINPUT110), .ZN(n664) );
  XNOR2_X2 U405 ( .A(n438), .B(n420), .ZN(n715) );
  XNOR2_X2 U406 ( .A(n374), .B(n373), .ZN(n438) );
  NOR2_X1 U407 ( .A1(G237), .A2(G953), .ZN(n433) );
  INV_X1 U408 ( .A(n528), .ZN(n558) );
  XNOR2_X1 U409 ( .A(n440), .B(G134), .ZN(n484) );
  XNOR2_X1 U410 ( .A(n363), .B(n362), .ZN(n452) );
  INV_X1 U411 ( .A(KEYINPUT92), .ZN(n362) );
  NOR2_X1 U412 ( .A1(n552), .A2(n361), .ZN(n403) );
  AND2_X1 U413 ( .A1(n550), .A2(n549), .ZN(n361) );
  AND2_X1 U414 ( .A1(n397), .A2(n394), .ZN(n393) );
  XNOR2_X1 U415 ( .A(G101), .B(G104), .ZN(n417) );
  INV_X1 U416 ( .A(G128), .ZN(n421) );
  NOR2_X1 U417 ( .A1(G902), .A2(n711), .ZN(n473) );
  XNOR2_X1 U418 ( .A(n726), .B(n442), .ZN(n615) );
  XOR2_X1 U419 ( .A(G125), .B(G140), .Z(n461) );
  INV_X1 U420 ( .A(KEYINPUT93), .ZN(n457) );
  XNOR2_X1 U421 ( .A(G116), .B(G107), .ZN(n477) );
  XOR2_X1 U422 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n479) );
  XNOR2_X1 U423 ( .A(n488), .B(n489), .ZN(n406) );
  XNOR2_X1 U424 ( .A(n561), .B(n560), .ZN(n685) );
  XNOR2_X1 U425 ( .A(n555), .B(n367), .ZN(n573) );
  INV_X1 U426 ( .A(KEYINPUT39), .ZN(n367) );
  INV_X1 U427 ( .A(KEYINPUT34), .ZN(n520) );
  NOR2_X1 U428 ( .A1(n656), .A2(n540), .ZN(n542) );
  NOR2_X1 U429 ( .A1(n706), .A2(G902), .ZN(n356) );
  BUF_X1 U430 ( .A(n656), .Z(n370) );
  AND2_X1 U431 ( .A1(n381), .A2(n384), .ZN(n360) );
  AND2_X1 U432 ( .A1(n379), .A2(n378), .ZN(n377) );
  OR2_X1 U433 ( .A1(n591), .A2(KEYINPUT96), .ZN(n378) );
  AND2_X1 U434 ( .A1(n617), .A2(G953), .ZN(n713) );
  XOR2_X1 U435 ( .A(KEYINPUT100), .B(n529), .Z(n665) );
  XNOR2_X1 U436 ( .A(G101), .B(KEYINPUT5), .ZN(n434) );
  XNOR2_X1 U437 ( .A(n419), .B(G119), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n375), .B(n376), .ZN(n374) );
  INV_X1 U439 ( .A(KEYINPUT72), .ZN(n419) );
  XOR2_X1 U440 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n426) );
  XNOR2_X1 U441 ( .A(KEYINPUT4), .B(G146), .ZN(n425) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n449) );
  AND2_X1 U443 ( .A1(n601), .A2(n366), .ZN(n475) );
  INV_X1 U444 ( .A(n540), .ZN(n366) );
  AND2_X1 U445 ( .A1(n591), .A2(KEYINPUT96), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n412), .B(KEYINPUT91), .ZN(n411) );
  INV_X1 U447 ( .A(KEYINPUT79), .ZN(n412) );
  XNOR2_X1 U448 ( .A(KEYINPUT16), .B(G122), .ZN(n420) );
  XNOR2_X1 U449 ( .A(KEYINPUT4), .B(G137), .ZN(n439) );
  AND2_X1 U450 ( .A1(n652), .A2(n533), .ZN(n534) );
  XNOR2_X1 U451 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n508) );
  INV_X1 U452 ( .A(KEYINPUT1), .ZN(n369) );
  INV_X1 U453 ( .A(KEYINPUT22), .ZN(n364) );
  AND2_X1 U454 ( .A1(n670), .A2(n577), .ZN(n578) );
  INV_X1 U455 ( .A(n516), .ZN(n600) );
  XNOR2_X1 U456 ( .A(n467), .B(n466), .ZN(n711) );
  XNOR2_X1 U457 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U458 ( .A(n484), .B(n483), .Z(n706) );
  XNOR2_X1 U459 ( .A(n352), .B(n487), .ZN(n404) );
  BUF_X1 U460 ( .A(n695), .Z(n709) );
  XNOR2_X1 U461 ( .A(n563), .B(n408), .ZN(n407) );
  OR2_X2 U462 ( .A1(n685), .A2(n562), .ZN(n409) );
  INV_X1 U463 ( .A(KEYINPUT111), .ZN(n408) );
  AND2_X1 U464 ( .A1(n556), .A2(n573), .ZN(n557) );
  XNOR2_X1 U465 ( .A(n556), .B(n495), .ZN(n638) );
  INV_X1 U466 ( .A(KEYINPUT105), .ZN(n495) );
  INV_X1 U467 ( .A(KEYINPUT97), .ZN(n593) );
  INV_X1 U468 ( .A(n713), .ZN(n357) );
  OR2_X1 U469 ( .A1(n513), .A2(n514), .ZN(n346) );
  OR2_X1 U470 ( .A1(n390), .A2(KEYINPUT0), .ZN(n347) );
  AND2_X1 U471 ( .A1(n358), .A2(n357), .ZN(n348) );
  AND2_X1 U472 ( .A1(n652), .A2(n399), .ZN(n349) );
  OR2_X1 U473 ( .A1(n516), .A2(n399), .ZN(n350) );
  INV_X1 U474 ( .A(n513), .ZN(n390) );
  XOR2_X1 U475 ( .A(KEYINPUT108), .B(n569), .Z(n351) );
  AND2_X1 U476 ( .A1(G214), .A2(n491), .ZN(n352) );
  AND2_X1 U477 ( .A1(n516), .A2(n652), .ZN(n353) );
  INV_X1 U478 ( .A(KEYINPUT96), .ZN(n389) );
  INV_X1 U479 ( .A(KEYINPUT102), .ZN(n399) );
  XNOR2_X1 U480 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n354) );
  XNOR2_X1 U481 ( .A(KEYINPUT62), .B(n615), .ZN(n355) );
  NAND2_X1 U482 ( .A1(n372), .A2(n609), .ZN(n687) );
  XNOR2_X1 U483 ( .A(n481), .B(n482), .ZN(n483) );
  NAND2_X1 U484 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U485 ( .A1(n592), .A2(n370), .ZN(n594) );
  NOR2_X1 U486 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U487 ( .A(n359), .B(n589), .ZN(n607) );
  NAND2_X1 U488 ( .A1(n596), .A2(n578), .ZN(n365) );
  XNOR2_X1 U489 ( .A(n616), .B(n355), .ZN(n358) );
  NAND2_X1 U490 ( .A1(n587), .A2(n588), .ZN(n359) );
  NAND2_X1 U491 ( .A1(n385), .A2(n387), .ZN(n384) );
  NAND2_X1 U492 ( .A1(n360), .A2(n377), .ZN(n592) );
  INV_X1 U493 ( .A(n387), .ZN(n383) );
  NOR2_X2 U494 ( .A1(n734), .A2(n735), .ZN(n564) );
  XNOR2_X2 U495 ( .A(n409), .B(n407), .ZN(n734) );
  NAND2_X1 U496 ( .A1(n553), .A2(n530), .ZN(n509) );
  XNOR2_X2 U497 ( .A(n368), .B(n432), .ZN(n553) );
  NAND2_X1 U498 ( .A1(n451), .A2(G902), .ZN(n363) );
  NOR2_X2 U499 ( .A1(n545), .A2(n562), .ZN(n639) );
  XNOR2_X1 U500 ( .A(n430), .B(n504), .ZN(n696) );
  XNOR2_X2 U501 ( .A(n365), .B(n364), .ZN(n584) );
  XNOR2_X2 U502 ( .A(n656), .B(KEYINPUT6), .ZN(n601) );
  NAND2_X1 U503 ( .A1(n545), .A2(n514), .ZN(n388) );
  NAND2_X1 U504 ( .A1(n696), .A2(n610), .ZN(n368) );
  NAND2_X1 U505 ( .A1(n349), .A2(n516), .ZN(n397) );
  XNOR2_X2 U506 ( .A(n543), .B(n369), .ZN(n516) );
  NAND2_X1 U507 ( .A1(n551), .A2(n403), .ZN(n402) );
  NAND2_X1 U508 ( .A1(n506), .A2(n341), .ZN(n551) );
  NAND2_X1 U509 ( .A1(n674), .A2(n596), .ZN(n521) );
  XNOR2_X1 U510 ( .A(n371), .B(n700), .ZN(G51) );
  NOR2_X2 U511 ( .A1(n699), .A2(n713), .ZN(n371) );
  NAND2_X1 U512 ( .A1(n396), .A2(KEYINPUT102), .ZN(n395) );
  AND2_X1 U513 ( .A1(n395), .A2(n601), .ZN(n394) );
  AND2_X1 U514 ( .A1(n372), .A2(n391), .ZN(n718) );
  NAND2_X1 U515 ( .A1(n380), .A2(n382), .ZN(n379) );
  INV_X1 U516 ( .A(n386), .ZN(n380) );
  NAND2_X1 U517 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U518 ( .A1(n528), .A2(n559), .ZN(n494) );
  XNOR2_X2 U519 ( .A(n583), .B(KEYINPUT32), .ZN(n736) );
  INV_X1 U520 ( .A(n652), .ZN(n396) );
  XNOR2_X2 U521 ( .A(n400), .B(n505), .ZN(n543) );
  XNOR2_X1 U522 ( .A(n402), .B(KEYINPUT69), .ZN(n566) );
  XNOR2_X1 U523 ( .A(n553), .B(KEYINPUT38), .ZN(n667) );
  INV_X1 U524 ( .A(n638), .ZN(n641) );
  NOR2_X1 U525 ( .A1(n341), .A2(n586), .ZN(n415) );
  XNOR2_X1 U526 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n416) );
  INV_X1 U527 ( .A(n650), .ZN(n577) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n567) );
  XNOR2_X1 U529 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U530 ( .A(n568), .B(n567), .ZN(n576) );
  XNOR2_X1 U531 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U532 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U534 ( .A(KEYINPUT42), .ZN(n563) );
  XNOR2_X1 U535 ( .A(n521), .B(n520), .ZN(n525) );
  XNOR2_X1 U536 ( .A(n431), .B(KEYINPUT85), .ZN(n432) );
  XNOR2_X1 U537 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U538 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  INV_X1 U539 ( .A(KEYINPUT75), .ZN(n418) );
  NAND2_X1 U540 ( .A1(G224), .A2(n391), .ZN(n423) );
  XNOR2_X1 U541 ( .A(n423), .B(G125), .ZN(n424) );
  XNOR2_X1 U542 ( .A(n440), .B(n424), .ZN(n428) );
  XNOR2_X1 U543 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U544 ( .A(n715), .B(n429), .ZN(n430) );
  OR2_X1 U545 ( .A1(G237), .A2(G902), .ZN(n498) );
  NAND2_X1 U546 ( .A1(n498), .A2(G210), .ZN(n431) );
  INV_X1 U547 ( .A(n553), .ZN(n571) );
  XNOR2_X1 U548 ( .A(n433), .B(KEYINPUT80), .ZN(n491) );
  NAND2_X1 U549 ( .A1(G210), .A2(n491), .ZN(n436) );
  XNOR2_X1 U550 ( .A(n434), .B(KEYINPUT78), .ZN(n435) );
  XNOR2_X1 U551 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U552 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U553 ( .A(n488), .B(n439), .ZN(n441) );
  XNOR2_X2 U554 ( .A(n484), .B(n441), .ZN(n726) );
  INV_X1 U555 ( .A(G902), .ZN(n443) );
  NAND2_X1 U556 ( .A1(n615), .A2(n443), .ZN(n445) );
  XOR2_X1 U557 ( .A(G472), .B(KEYINPUT76), .Z(n444) );
  XNOR2_X2 U558 ( .A(n445), .B(n444), .ZN(n656) );
  XOR2_X1 U559 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n448) );
  NAND2_X1 U560 ( .A1(G234), .A2(n610), .ZN(n446) );
  XNOR2_X1 U561 ( .A(KEYINPUT20), .B(n446), .ZN(n468) );
  NAND2_X1 U562 ( .A1(n468), .A2(G221), .ZN(n447) );
  XNOR2_X1 U563 ( .A(n448), .B(n447), .ZN(n650) );
  XOR2_X1 U564 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n450) );
  XNOR2_X1 U565 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U566 ( .A1(G952), .A2(n451), .ZN(n682) );
  NOR2_X1 U567 ( .A1(G953), .A2(n682), .ZN(n512) );
  NAND2_X1 U568 ( .A1(G953), .A2(n452), .ZN(n510) );
  NOR2_X1 U569 ( .A1(G900), .A2(n510), .ZN(n453) );
  NOR2_X1 U570 ( .A1(n512), .A2(n453), .ZN(n532) );
  NOR2_X1 U571 ( .A1(n650), .A2(n532), .ZN(n454) );
  XNOR2_X1 U572 ( .A(n454), .B(KEYINPUT70), .ZN(n474) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(G137), .Z(n456) );
  XNOR2_X1 U574 ( .A(G146), .B(G128), .ZN(n455) );
  XNOR2_X1 U575 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U576 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U577 ( .A(n462), .B(n727), .ZN(n467) );
  NAND2_X1 U578 ( .A1(G234), .A2(n391), .ZN(n463) );
  XOR2_X1 U579 ( .A(KEYINPUT8), .B(n463), .Z(n476) );
  NAND2_X1 U580 ( .A1(n476), .A2(G221), .ZN(n465) );
  XNOR2_X1 U581 ( .A(KEYINPUT74), .B(KEYINPUT24), .ZN(n464) );
  NAND2_X1 U582 ( .A1(n468), .A2(G217), .ZN(n471) );
  XNOR2_X1 U583 ( .A(KEYINPUT94), .B(KEYINPUT81), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n469), .B(KEYINPUT25), .ZN(n470) );
  NAND2_X1 U585 ( .A1(n474), .A2(n649), .ZN(n540) );
  XNOR2_X1 U586 ( .A(n475), .B(KEYINPUT106), .ZN(n496) );
  NAND2_X1 U587 ( .A1(G217), .A2(n476), .ZN(n482) );
  XOR2_X1 U588 ( .A(KEYINPUT9), .B(G122), .Z(n478) );
  XNOR2_X1 U589 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U590 ( .A(KEYINPUT13), .B(G475), .ZN(n493) );
  INV_X1 U591 ( .A(n727), .ZN(n490) );
  XOR2_X1 U592 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n489) );
  XOR2_X1 U593 ( .A(G122), .B(G104), .Z(n486) );
  XNOR2_X1 U594 ( .A(G113), .B(G143), .ZN(n485) );
  XNOR2_X1 U595 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U596 ( .A1(G902), .A2(n701), .ZN(n492) );
  XNOR2_X1 U597 ( .A(n493), .B(n492), .ZN(n559) );
  NAND2_X1 U598 ( .A1(n496), .A2(n638), .ZN(n497) );
  NAND2_X1 U599 ( .A1(G214), .A2(n498), .ZN(n530) );
  NAND2_X1 U600 ( .A1(n499), .A2(n530), .ZN(n569) );
  XNOR2_X1 U601 ( .A(n500), .B(KEYINPUT36), .ZN(n506) );
  NAND2_X1 U602 ( .A1(n391), .A2(G227), .ZN(n502) );
  XNOR2_X1 U603 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U604 ( .A(KEYINPUT71), .B(G469), .ZN(n505) );
  XOR2_X1 U605 ( .A(G125), .B(KEYINPUT37), .Z(n507) );
  XNOR2_X1 U606 ( .A(n551), .B(n507), .ZN(G27) );
  XNOR2_X2 U607 ( .A(n509), .B(n508), .ZN(n545) );
  NOR2_X1 U608 ( .A1(G898), .A2(n510), .ZN(n511) );
  NOR2_X1 U609 ( .A1(n512), .A2(n511), .ZN(n513) );
  INV_X1 U610 ( .A(KEYINPUT0), .ZN(n514) );
  NOR2_X1 U611 ( .A1(n649), .A2(n650), .ZN(n515) );
  XNOR2_X2 U612 ( .A(n515), .B(KEYINPUT66), .ZN(n652) );
  XNOR2_X1 U613 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n518) );
  INV_X1 U614 ( .A(KEYINPUT90), .ZN(n517) );
  XNOR2_X1 U615 ( .A(n518), .B(n517), .ZN(n519) );
  AND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n523) );
  INV_X1 U617 ( .A(KEYINPUT104), .ZN(n522) );
  XNOR2_X1 U618 ( .A(n523), .B(n522), .ZN(n536) );
  INV_X1 U619 ( .A(n536), .ZN(n524) );
  XNOR2_X1 U620 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n526) );
  XNOR2_X1 U621 ( .A(n588), .B(G122), .ZN(G24) );
  NOR2_X1 U622 ( .A1(n559), .A2(n528), .ZN(n633) );
  NOR2_X1 U623 ( .A1(n556), .A2(n633), .ZN(n529) );
  INV_X1 U624 ( .A(n665), .ZN(n548) );
  NAND2_X1 U625 ( .A1(n548), .A2(KEYINPUT47), .ZN(n538) );
  INV_X1 U626 ( .A(n530), .ZN(n668) );
  OR2_X1 U627 ( .A1(n668), .A2(n656), .ZN(n531) );
  XOR2_X1 U628 ( .A(KEYINPUT30), .B(n531), .Z(n535) );
  NOR2_X1 U629 ( .A1(n543), .A2(n532), .ZN(n533) );
  NAND2_X1 U630 ( .A1(n535), .A2(n534), .ZN(n554) );
  NOR2_X1 U631 ( .A1(n536), .A2(n554), .ZN(n537) );
  NAND2_X1 U632 ( .A1(n345), .A2(n537), .ZN(n637) );
  NAND2_X1 U633 ( .A1(n538), .A2(n637), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n539), .B(KEYINPUT86), .ZN(n552) );
  INV_X1 U635 ( .A(KEYINPUT67), .ZN(n546) );
  XOR2_X1 U636 ( .A(KEYINPUT28), .B(KEYINPUT109), .Z(n541) );
  XNOR2_X1 U637 ( .A(n542), .B(n541), .ZN(n544) );
  INV_X1 U638 ( .A(n543), .ZN(n590) );
  NAND2_X1 U639 ( .A1(n544), .A2(n590), .ZN(n562) );
  NAND2_X1 U640 ( .A1(n546), .A2(n639), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n547), .B(KEYINPUT47), .ZN(n550) );
  NAND2_X1 U642 ( .A1(n548), .A2(n639), .ZN(n549) );
  NOR2_X1 U643 ( .A1(n554), .A2(n667), .ZN(n555) );
  XNOR2_X1 U644 ( .A(n557), .B(KEYINPUT40), .ZN(n735) );
  NOR2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n670) );
  NAND2_X1 U646 ( .A1(n664), .A2(n670), .ZN(n561) );
  INV_X1 U647 ( .A(KEYINPUT41), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n564), .B(KEYINPUT46), .ZN(n565) );
  NAND2_X1 U649 ( .A1(n565), .A2(n566), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n351), .A2(n600), .ZN(n570) );
  XNOR2_X1 U651 ( .A(n570), .B(KEYINPUT43), .ZN(n572) );
  AND2_X1 U652 ( .A1(n572), .A2(n571), .ZN(n648) );
  INV_X1 U653 ( .A(n648), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n573), .A2(n633), .ZN(n646) );
  AND2_X1 U655 ( .A1(n574), .A2(n646), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n576), .A2(n575), .ZN(n725) );
  INV_X1 U657 ( .A(n725), .ZN(n609) );
  XNOR2_X1 U658 ( .A(KEYINPUT83), .B(n601), .ZN(n579) );
  NAND2_X1 U659 ( .A1(n579), .A2(n649), .ZN(n580) );
  NOR2_X1 U660 ( .A1(n580), .A2(n600), .ZN(n581) );
  XNOR2_X1 U661 ( .A(n581), .B(KEYINPUT82), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n584), .A2(n582), .ZN(n583) );
  INV_X1 U663 ( .A(n370), .ZN(n595) );
  INV_X1 U664 ( .A(n649), .ZN(n585) );
  OR2_X1 U665 ( .A1(n595), .A2(n585), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n584), .A2(n415), .ZN(n632) );
  INV_X1 U667 ( .A(KEYINPUT44), .ZN(n589) );
  AND2_X1 U668 ( .A1(n652), .A2(n590), .ZN(n591) );
  AND2_X1 U669 ( .A1(n353), .A2(n595), .ZN(n659) );
  NAND2_X1 U670 ( .A1(n596), .A2(n659), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT31), .B(n597), .Z(n643) );
  NAND2_X1 U672 ( .A1(n629), .A2(n643), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n598), .A2(n665), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT101), .ZN(n605) );
  AND2_X1 U675 ( .A1(n584), .A2(n600), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n601), .A2(n649), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n624) );
  INV_X1 U678 ( .A(n624), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n687), .B(KEYINPUT2), .ZN(n612) );
  INV_X1 U680 ( .A(n610), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U682 ( .A(KEYINPUT64), .ZN(n613) );
  XNOR2_X2 U683 ( .A(n614), .B(n613), .ZN(n695) );
  NAND2_X1 U684 ( .A1(n695), .A2(G472), .ZN(n616) );
  INV_X1 U685 ( .A(G952), .ZN(n617) );
  XOR2_X1 U686 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n618) );
  XNOR2_X1 U687 ( .A(n348), .B(n618), .ZN(G57) );
  NAND2_X1 U688 ( .A1(n709), .A2(G469), .ZN(n622) );
  XOR2_X1 U689 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U692 ( .A1(n623), .A2(n713), .ZN(G54) );
  XNOR2_X1 U693 ( .A(G101), .B(n624), .ZN(G3) );
  NOR2_X1 U694 ( .A1(n641), .A2(n629), .ZN(n626) );
  XNOR2_X1 U695 ( .A(G104), .B(KEYINPUT113), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n626), .B(n625), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n628) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT27), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n631) );
  INV_X1 U700 ( .A(n633), .ZN(n644) );
  NOR2_X1 U701 ( .A1(n644), .A2(n629), .ZN(n630) );
  XOR2_X1 U702 ( .A(n631), .B(n630), .Z(G9) );
  XNOR2_X1 U703 ( .A(G110), .B(n632), .ZN(G12) );
  XOR2_X1 U704 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n635) );
  NAND2_X1 U705 ( .A1(n639), .A2(n633), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  XOR2_X1 U707 ( .A(G128), .B(n636), .Z(G30) );
  XNOR2_X1 U708 ( .A(G143), .B(n637), .ZN(G45) );
  NAND2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(G146), .ZN(G48) );
  NOR2_X1 U711 ( .A1(n641), .A2(n643), .ZN(n642) );
  XOR2_X1 U712 ( .A(G113), .B(n642), .Z(G15) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U714 ( .A(G116), .B(n645), .Z(G18) );
  XNOR2_X1 U715 ( .A(G134), .B(KEYINPUT116), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G36) );
  XOR2_X1 U717 ( .A(G140), .B(n648), .Z(G42) );
  NAND2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT49), .B(n651), .ZN(n658) );
  NOR2_X1 U720 ( .A1(n652), .A2(n341), .ZN(n654) );
  XNOR2_X1 U721 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U723 ( .A1(n370), .A2(n655), .ZN(n657) );
  NOR2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n660) );
  NOR2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U726 ( .A(n661), .B(KEYINPUT51), .Z(n662) );
  XNOR2_X1 U727 ( .A(KEYINPUT118), .B(n662), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n685), .A2(n663), .ZN(n678) );
  NAND2_X1 U729 ( .A1(n665), .A2(n344), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT119), .B(n666), .Z(n672) );
  NAND2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U734 ( .A(KEYINPUT120), .B(n673), .Z(n675) );
  INV_X1 U735 ( .A(n674), .ZN(n684) );
  NOR2_X1 U736 ( .A1(n675), .A2(n684), .ZN(n676) );
  XOR2_X1 U737 ( .A(n676), .B(KEYINPUT121), .Z(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U739 ( .A(KEYINPUT52), .B(n679), .Z(n680) );
  XOR2_X1 U740 ( .A(KEYINPUT122), .B(n680), .Z(n681) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U742 ( .A(KEYINPUT123), .B(n683), .Z(n692) );
  NOR2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n686), .A2(G953), .ZN(n690) );
  NOR2_X1 U745 ( .A1(n343), .A2(KEYINPUT87), .ZN(n688) );
  XOR2_X1 U746 ( .A(n688), .B(KEYINPUT2), .Z(n689) );
  NAND2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U749 ( .A(KEYINPUT53), .B(KEYINPUT124), .ZN(n693) );
  XNOR2_X1 U750 ( .A(n694), .B(n693), .ZN(G75) );
  NAND2_X1 U751 ( .A1(n695), .A2(G210), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n696), .B(n416), .ZN(n697) );
  XOR2_X1 U753 ( .A(KEYINPUT56), .B(KEYINPUT125), .Z(n700) );
  NAND2_X1 U754 ( .A1(n695), .A2(G475), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X2 U756 ( .A1(n704), .A2(n713), .ZN(n705) );
  XNOR2_X1 U757 ( .A(n705), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U758 ( .A1(n709), .A2(G478), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n713), .A2(n708), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n709), .A2(G217), .ZN(n710) );
  XNOR2_X1 U762 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n713), .A2(n712), .ZN(G66) );
  NOR2_X1 U764 ( .A1(G898), .A2(n391), .ZN(n717) );
  XOR2_X1 U765 ( .A(n714), .B(n715), .Z(n716) );
  NOR2_X1 U766 ( .A1(n717), .A2(n716), .ZN(n724) );
  XOR2_X1 U767 ( .A(n718), .B(KEYINPUT126), .Z(n722) );
  NAND2_X1 U768 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n720), .A2(G898), .ZN(n721) );
  NAND2_X1 U771 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(G69) );
  XOR2_X1 U773 ( .A(n727), .B(n726), .Z(n729) );
  XNOR2_X1 U774 ( .A(n725), .B(n729), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(n391), .ZN(n733) );
  XNOR2_X1 U776 ( .A(n729), .B(G227), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U779 ( .A1(n733), .A2(n732), .ZN(G72) );
  XOR2_X1 U780 ( .A(n734), .B(G137), .Z(G39) );
  XOR2_X1 U781 ( .A(G131), .B(n735), .Z(G33) );
  XNOR2_X1 U782 ( .A(n736), .B(G119), .ZN(G21) );
endmodule

