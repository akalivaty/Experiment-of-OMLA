//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(KEYINPUT93), .B2(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n189), .B1(KEYINPUT93), .B2(new_n188), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT9), .B(G234), .ZN(new_n191));
  INV_X1    g005(.A(G217), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n191), .A2(new_n192), .A3(G953), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT64), .A2(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT64), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n202), .B2(G128), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR4_X1   g018(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT92), .A4(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n195), .B(new_n198), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G122), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G122), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT76), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n211), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n206), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT13), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n203), .B2(new_n205), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT64), .B(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT92), .B1(new_n221), .B2(new_n204), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n202), .A2(new_n199), .A3(G128), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT13), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n224), .A3(new_n198), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n218), .B1(G134), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n211), .A2(new_n216), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n209), .A2(KEYINPUT14), .A3(G122), .ZN(new_n228));
  OAI211_X1 g042(.A(G107), .B(new_n228), .C1(new_n211), .C2(KEYINPUT14), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n223), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n198), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G134), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(new_n233), .B2(new_n206), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n194), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n230), .ZN(new_n236));
  INV_X1    g050(.A(new_n206), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n195), .B1(new_n231), .B2(new_n198), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n197), .B1(new_n231), .B2(new_n219), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n195), .B1(new_n240), .B2(new_n224), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n239), .B(new_n193), .C1(new_n241), .C2(new_n218), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G902), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT94), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT94), .ZN(new_n246));
  AOI211_X1 g060(.A(new_n246), .B(G902), .C1(new_n235), .C2(new_n242), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n190), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n190), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n235), .B2(new_n242), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n251), .B2(new_n246), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT95), .ZN(new_n254));
  NAND2_X1  g068(.A1(G234), .A2(G237), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n255), .A2(G952), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n255), .A2(G902), .A3(G953), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT21), .B(G898), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT95), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n248), .A2(new_n262), .A3(new_n252), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n254), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(G475), .A2(G902), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G113), .B(G122), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT89), .B(G104), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n267), .B(new_n268), .Z(new_n269));
  XNOR2_X1  g083(.A(G125), .B(G140), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT72), .A2(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT72), .A2(G125), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(G140), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n276));
  INV_X1    g090(.A(G125), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G140), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n273), .A2(KEYINPUT73), .A3(G140), .A4(new_n274), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n272), .B1(new_n282), .B2(new_n271), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT18), .A2(G131), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(KEYINPUT86), .ZN(new_n286));
  INV_X1    g100(.A(G237), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n256), .A3(G214), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT64), .A2(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT64), .A2(G143), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(G143), .A2(G214), .ZN(new_n292));
  NOR4_X1   g106(.A1(new_n292), .A2(KEYINPUT85), .A3(G237), .A4(G953), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n294));
  AND2_X1   g108(.A1(G143), .A2(G214), .ZN(new_n295));
  NOR2_X1   g109(.A1(G237), .A2(G953), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n291), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n285), .A2(new_n284), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n283), .B(new_n300), .C1(new_n286), .C2(new_n298), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n287), .A2(new_n256), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT85), .B1(new_n303), .B2(new_n292), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n295), .A2(new_n296), .A3(new_n294), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n304), .A2(new_n305), .B1(new_n202), .B2(new_n288), .ZN(new_n306));
  INV_X1    g120(.A(G131), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT17), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n298), .A2(KEYINPUT88), .A3(G131), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n307), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT90), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n280), .B2(new_n281), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT72), .A2(G125), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT72), .A2(G125), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n319), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n271), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n278), .B1(new_n319), .B2(G140), .ZN(new_n322));
  INV_X1    g136(.A(new_n281), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT16), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n320), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(G146), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n308), .A2(new_n310), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT17), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n314), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n312), .A2(new_n313), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n269), .B(new_n301), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n307), .B2(new_n306), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT19), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n270), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n282), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n326), .B1(new_n336), .B2(G146), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n301), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n269), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n266), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT91), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n341), .A2(new_n342), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n332), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n312), .A2(new_n313), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n327), .A3(new_n314), .A4(new_n329), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n269), .B1(new_n351), .B2(new_n301), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n244), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G475), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n264), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G214), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT2), .B(G113), .Z(new_n359));
  XNOR2_X1  g173(.A(G116), .B(G119), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n360), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n212), .B1(new_n365), .B2(G104), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(KEYINPUT3), .B2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n213), .A2(new_n215), .A3(new_n365), .A4(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G101), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n375));
  AND4_X1   g189(.A1(KEYINPUT77), .A2(new_n370), .A3(new_n375), .A4(G101), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n368), .B2(new_n369), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT77), .B1(new_n377), .B2(new_n375), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n364), .B(new_n374), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n370), .A2(new_n375), .A3(G101), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(KEYINPUT77), .A3(new_n375), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(KEYINPUT80), .A3(new_n364), .A4(new_n374), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n360), .A2(KEYINPUT5), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n209), .A2(KEYINPUT5), .A3(G119), .ZN(new_n390));
  INV_X1    g204(.A(G113), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n372), .B1(G104), .B2(G107), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n216), .B2(G104), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n373), .A2(new_n393), .A3(new_n361), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT81), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n397), .B1(new_n381), .B2(new_n387), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n400), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n271), .A2(G143), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n202), .B2(G146), .ZN(new_n409));
  AND2_X1   g223(.A1(KEYINPUT0), .A2(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n271), .B1(new_n200), .B2(new_n201), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n196), .A2(G146), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(KEYINPUT0), .A2(G128), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n318), .B2(new_n317), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n289), .A2(G146), .A3(new_n290), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n407), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n407), .A2(KEYINPUT1), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n412), .A2(new_n413), .B1(new_n424), .B2(G128), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n319), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G224), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(G953), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n427), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n399), .A2(new_n403), .A3(new_n401), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n406), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n373), .A2(new_n395), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n389), .B(KEYINPUT82), .Z(new_n435));
  XOR2_X1   g249(.A(new_n392), .B(KEYINPUT83), .Z(new_n436));
  OAI21_X1  g250(.A(new_n361), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n434), .B1(new_n437), .B2(KEYINPUT84), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(KEYINPUT84), .B2(new_n437), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n400), .B(KEYINPUT8), .Z(new_n440));
  AND2_X1   g254(.A1(new_n393), .A2(new_n361), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n434), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n419), .A2(KEYINPUT7), .A3(new_n430), .A4(new_n426), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n427), .B1(new_n444), .B2(new_n429), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n439), .A2(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n404), .A2(new_n400), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n433), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n433), .A2(new_n448), .A3(new_n450), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n358), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G221), .B1(new_n191), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G469), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n244), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G140), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n256), .A2(G227), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n459), .B(new_n460), .Z(new_n461));
  OAI211_X1 g275(.A(new_n418), .B(new_n374), .C1(new_n376), .C2(new_n378), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n373), .A2(new_n395), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n204), .B1(new_n412), .B2(KEYINPUT1), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n422), .B1(new_n464), .B2(new_n409), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT11), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n195), .B2(G137), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n195), .A2(G137), .ZN(new_n471));
  INV_X1    g285(.A(G137), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT11), .A3(G134), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G131), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n470), .A2(new_n473), .A3(new_n307), .A4(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  INV_X1    g293(.A(new_n425), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n422), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n463), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n462), .A2(new_n468), .A3(new_n478), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n466), .A2(new_n467), .B1(new_n481), .B2(new_n463), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n478), .B1(new_n485), .B2(new_n462), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n461), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n461), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n434), .A2(new_n422), .A3(new_n480), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n466), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n490), .A2(KEYINPUT12), .A3(new_n477), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n490), .B2(new_n477), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n488), .B(new_n483), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n458), .B1(new_n494), .B2(new_n457), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n483), .A2(new_n488), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT79), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT79), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n483), .A2(new_n498), .A3(new_n488), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n462), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n477), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n491), .A2(new_n492), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n461), .B1(new_n503), .B2(new_n484), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(G469), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n456), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n356), .A2(KEYINPUT96), .A3(new_n454), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n248), .A2(new_n262), .A3(new_n252), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n262), .B1(new_n248), .B2(new_n252), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n509), .A2(new_n510), .A3(new_n260), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n353), .A2(G475), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n345), .B1(new_n341), .B2(new_n342), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n341), .A2(new_n342), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n515), .B2(new_n346), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n433), .A2(new_n448), .A3(new_n450), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n450), .B1(new_n433), .B2(new_n448), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n506), .B(new_n357), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n508), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n321), .A2(new_n326), .ZN(new_n522));
  XOR2_X1   g336(.A(G119), .B(G128), .Z(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT24), .B(G110), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT71), .B1(new_n526), .B2(G128), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n527), .A2(KEYINPUT23), .B1(new_n526), .B2(G128), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(KEYINPUT23), .B2(new_n527), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n525), .B1(new_n529), .B2(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n524), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT74), .B(G110), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n532), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n326), .A2(new_n272), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n256), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT75), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT22), .B(G137), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n531), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n531), .B2(new_n535), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n192), .B1(G234), .B2(new_n244), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n542), .B2(G902), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT25), .B(new_n244), .C1(new_n540), .C2(new_n541), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n550), .B2(new_n543), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(G472), .A2(G902), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n477), .A2(new_n411), .A3(new_n417), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n472), .A2(G134), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n195), .A2(G137), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n476), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n423), .B2(new_n425), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n362), .A2(new_n363), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n554), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT28), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT68), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT26), .B(G101), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n296), .A2(G210), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT67), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT67), .ZN(new_n577));
  INV_X1    g391(.A(new_n574), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n573), .A2(new_n578), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n570), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT65), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT30), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n585), .B(new_n586), .C1(new_n554), .C2(new_n559), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g402(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n554), .A2(new_n559), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n364), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT31), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n564), .A4(new_n575), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n554), .A2(new_n559), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT65), .A3(KEYINPUT30), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n590), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n561), .B1(new_n598), .B2(new_n364), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n599), .B2(new_n575), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n553), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT32), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT32), .B(new_n553), .C1(new_n595), .C2(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G472), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n575), .A2(KEYINPUT29), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n244), .B1(new_n570), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n575), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n560), .B1(new_n597), .B2(new_n590), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n561), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT29), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n563), .A2(new_n567), .A3(new_n582), .A4(new_n569), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT69), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n608), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT69), .A4(new_n612), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n606), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT70), .B1(new_n605), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n616), .A2(new_n617), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT70), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n603), .A4(new_n604), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n552), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n507), .A2(new_n521), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  OR3_X1    g441(.A1(new_n243), .A2(new_n627), .A3(KEYINPUT33), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(KEYINPUT33), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n243), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n187), .A2(G902), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n633), .A2(new_n634), .B1(new_n187), .B2(new_n251), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n348), .B2(new_n354), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n454), .A2(new_n636), .A3(new_n261), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n592), .A2(new_n564), .A3(new_n575), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT31), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n594), .A3(new_n584), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n244), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G472), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n506), .A2(new_n551), .A3(new_n601), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  OAI211_X1 g460(.A(new_n261), .B(new_n357), .C1(new_n518), .C2(new_n519), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n347), .A2(new_n343), .B1(new_n353), .B2(G475), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n510), .B2(new_n509), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n647), .A2(new_n643), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT35), .B(G107), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NAND2_X1  g466(.A1(new_n550), .A2(new_n543), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n531), .A2(new_n535), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n544), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n642), .A2(new_n601), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n507), .A2(new_n521), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n506), .A2(new_n658), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n619), .B2(new_n623), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n257), .B1(new_n258), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n648), .B(new_n669), .C1(new_n510), .C2(new_n509), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n666), .A2(new_n454), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n452), .A2(new_n453), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT38), .Z(new_n675));
  NOR2_X1   g489(.A1(new_n509), .A2(new_n510), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n516), .A2(new_n676), .A3(new_n358), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n604), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT32), .B1(new_n640), .B2(new_n553), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n561), .A2(new_n562), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n599), .A2(new_n575), .B1(new_n583), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n683), .B2(G902), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n658), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n675), .A2(new_n678), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n668), .B(KEYINPUT39), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n506), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT98), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n221), .ZN(G45));
  INV_X1    g508(.A(new_n635), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n341), .A2(new_n345), .A3(new_n342), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n513), .A3(new_n514), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n695), .B(new_n669), .C1(new_n697), .C2(new_n512), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT99), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT99), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n636), .A2(new_n700), .A3(new_n669), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n666), .A2(new_n699), .A3(new_n454), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(new_n355), .A2(new_n695), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n647), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n487), .A2(new_n493), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n457), .A3(new_n244), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n494), .A2(new_n457), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n456), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n624), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT100), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(G15));
  NOR2_X1   g528(.A1(new_n647), .A2(new_n649), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n624), .A2(new_n715), .A3(new_n710), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AOI21_X1  g531(.A(new_n622), .B1(new_n681), .B2(new_n621), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n605), .A2(KEYINPUT70), .A3(new_n618), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n658), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n454), .A2(new_n516), .A3(new_n511), .A4(new_n710), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT101), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n710), .B(new_n357), .C1(new_n518), .C2(new_n519), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n517), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n659), .B1(new_n619), .B2(new_n623), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n641), .B2(G472), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n731), .B(new_n606), .C1(new_n640), .C2(new_n244), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n601), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n640), .A2(KEYINPUT102), .A3(new_n553), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n733), .A2(new_n552), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n710), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n647), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n516), .A2(new_n676), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NOR3_X1   g557(.A1(new_n733), .A2(new_n659), .A3(new_n737), .ZN(new_n744));
  INV_X1    g558(.A(new_n723), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n699), .A3(new_n701), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n619), .A2(new_n623), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n452), .A2(new_n357), .A3(new_n453), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n458), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n505), .A2(new_n707), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n455), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n506), .A2(KEYINPUT104), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n749), .A2(new_n551), .A3(new_n751), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n699), .A2(new_n701), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n748), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n755), .B(new_n456), .C1(new_n495), .C2(new_n505), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT104), .B1(new_n753), .B2(new_n455), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n748), .A3(new_n750), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n604), .B(KEYINPUT105), .Z(new_n766));
  NOR2_X1   g580(.A1(new_n618), .A2(new_n680), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n552), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n701), .A3(new_n699), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT106), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n761), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n307), .ZN(G33));
  AOI21_X1  g589(.A(new_n750), .B1(new_n756), .B2(new_n757), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n624), .A2(new_n776), .A3(new_n671), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n195), .ZN(G36));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n779), .B(KEYINPUT43), .C1(new_n355), .C2(new_n635), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n516), .A2(new_n695), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n660), .A2(new_n658), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(KEYINPUT44), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(new_n783), .A3(new_n785), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n750), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n502), .A2(new_n504), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n457), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n504), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n752), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n708), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n456), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n786), .A2(new_n789), .A3(KEYINPUT108), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n792), .A2(new_n688), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NOR2_X1   g619(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n807), .B(new_n456), .C1(new_n800), .C2(new_n801), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n749), .A2(new_n551), .A3(new_n750), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n701), .A3(new_n699), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n806), .A2(new_n808), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n814), .B1(new_n815), .B2(new_n811), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NOR2_X1   g632(.A1(new_n708), .A2(new_n709), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT49), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n552), .A2(new_n358), .A3(new_n456), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n695), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n681), .A2(new_n684), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n516), .A3(new_n675), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n675), .A2(new_n358), .A3(new_n710), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n784), .A2(new_n257), .ZN(new_n829));
  INV_X1    g643(.A(new_n738), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(KEYINPUT50), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n551), .A2(new_n257), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n823), .A2(new_n750), .A3(new_n739), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n355), .A2(new_n695), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n784), .A2(new_n257), .A3(new_n710), .A4(new_n751), .ZN(new_n841));
  INV_X1    g655(.A(new_n744), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT116), .Z(new_n844));
  NOR3_X1   g658(.A1(new_n829), .A2(new_n830), .A3(new_n750), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n819), .A2(new_n456), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT114), .Z(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n809), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n836), .A2(new_n840), .A3(new_n844), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT48), .ZN(new_n852));
  INV_X1    g666(.A(new_n768), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n841), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n831), .A2(new_n745), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n852), .B1(new_n841), .B2(new_n853), .ZN(new_n856));
  INV_X1    g670(.A(G952), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n857), .B(G953), .C1(new_n838), .C2(new_n636), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n846), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n845), .B1(new_n809), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n844), .A2(KEYINPUT51), .A3(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n834), .A2(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n851), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n507), .B(new_n521), .C1(new_n624), .C2(new_n661), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n643), .B1(new_n637), .B2(KEYINPUT110), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n705), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n720), .A2(KEYINPUT101), .A3(new_n721), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n868), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n647), .A2(new_n643), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n253), .A2(KEYINPUT111), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n248), .A2(new_n878), .A3(new_n252), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n355), .A2(new_n880), .A3(KEYINPUT112), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n248), .A2(new_n878), .A3(new_n252), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n878), .B1(new_n248), .B2(new_n252), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n882), .B1(new_n516), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n876), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n711), .A2(new_n716), .A3(new_n742), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n875), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n880), .A2(new_n648), .A3(new_n669), .ZN(new_n890));
  INV_X1    g704(.A(new_n665), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n749), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n730), .ZN(new_n893));
  INV_X1    g707(.A(new_n732), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n737), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n758), .A3(new_n658), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n760), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n777), .B1(new_n897), .B2(new_n751), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n889), .A2(new_n771), .A3(new_n773), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n668), .B(KEYINPUT113), .Z(new_n900));
  NOR2_X1   g714(.A1(new_n754), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n677), .A2(new_n674), .A3(new_n685), .A4(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n702), .A2(new_n746), .A3(new_n672), .A4(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n867), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n722), .A2(new_n727), .B1(new_n871), .B2(new_n869), .ZN(new_n908));
  AND4_X1   g722(.A1(new_n711), .A2(new_n716), .A3(new_n742), .A4(new_n887), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n898), .A2(new_n908), .A3(new_n909), .A4(new_n868), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n774), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n746), .A2(new_n672), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT52), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n867), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n905), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n866), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n911), .B2(new_n905), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n770), .A2(new_n913), .A3(KEYINPUT53), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n905), .A2(new_n889), .A3(new_n918), .A4(new_n898), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n917), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n865), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(G952), .A2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n825), .B1(new_n922), .B2(new_n923), .ZN(G75));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n857), .A2(G953), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT118), .ZN(new_n927));
  INV_X1    g741(.A(G210), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n928), .B(new_n244), .C1(new_n907), .C2(new_n919), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n406), .A2(new_n432), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n431), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n927), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n932), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n907), .A2(new_n919), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(G210), .A3(G902), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n925), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n932), .B1(new_n929), .B2(KEYINPUT56), .ZN(new_n943));
  INV_X1    g757(.A(new_n927), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n939), .B2(new_n934), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n945), .A3(KEYINPUT119), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(new_n946), .ZN(G51));
  OAI21_X1  g761(.A(KEYINPUT54), .B1(new_n917), .B2(new_n920), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n907), .A2(new_n866), .A3(new_n919), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n938), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n458), .B(KEYINPUT57), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n706), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n917), .A2(new_n920), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n244), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n796), .A3(new_n795), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n944), .B1(new_n955), .B2(new_n958), .ZN(G54));
  NAND3_X1  g773(.A1(new_n957), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n332), .A2(new_n340), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n957), .A2(KEYINPUT58), .A3(G475), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n944), .B1(new_n962), .B2(new_n964), .ZN(G60));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT59), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n921), .B2(new_n916), .ZN(new_n969));
  INV_X1    g783(.A(new_n633), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n944), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n951), .A2(new_n633), .A3(new_n952), .A4(new_n968), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n542), .B1(new_n956), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n938), .A2(new_n656), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n927), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n976), .A2(KEYINPUT61), .A3(new_n927), .A4(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n259), .B2(new_n428), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n889), .B2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n930), .B1(G898), .B2(new_n256), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT121), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  AND2_X1   g802(.A1(new_n690), .A2(new_n751), .ZN(new_n989));
  OR3_X1    g803(.A1(new_n881), .A2(new_n886), .A3(new_n636), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n990), .A3(new_n624), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT122), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT122), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(new_n990), .A3(new_n993), .A4(new_n624), .ZN(new_n994));
  AOI22_X1  g808(.A1(new_n813), .A2(new_n816), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n693), .ZN(new_n996));
  INV_X1    g810(.A(new_n912), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n702), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT62), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n693), .A2(new_n1000), .A3(new_n702), .A4(new_n997), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n995), .A2(new_n999), .A3(new_n804), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n256), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n598), .B(new_n336), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n256), .A2(G900), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT123), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n802), .A2(new_n688), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n768), .A2(new_n674), .A3(new_n677), .ZN(new_n1009));
  OAI22_X1  g823(.A1(new_n1008), .A2(new_n1009), .B1(new_n670), .B2(new_n759), .ZN(new_n1010));
  AOI211_X1 g824(.A(new_n998), .B(new_n1010), .C1(new_n813), .C2(new_n816), .ZN(new_n1011));
  INV_X1    g825(.A(new_n774), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n804), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1007), .B1(new_n1013), .B2(new_n256), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1005), .B1(new_n1014), .B2(new_n1004), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n256), .B1(G227), .B2(G900), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G72));
  XNOR2_X1  g831(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n606), .A2(new_n244), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1018), .B(new_n1019), .Z(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n638), .B2(new_n611), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT127), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n907), .B2(new_n915), .ZN(new_n1024));
  INV_X1    g838(.A(new_n599), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n575), .ZN(new_n1026));
  INV_X1    g840(.A(new_n889), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1020), .B1(new_n1002), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT125), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g844(.A(KEYINPUT125), .B(new_n1020), .C1(new_n1002), .C2(new_n1027), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1011), .A2(new_n1012), .A3(new_n804), .A4(new_n889), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n1020), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1025), .A2(new_n575), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(KEYINPUT126), .A3(new_n927), .ZN(new_n1036));
  INV_X1    g850(.A(KEYINPUT126), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1034), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n1032), .B2(new_n1020), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1037), .B1(new_n1039), .B2(new_n944), .ZN(new_n1040));
  AOI221_X4 g854(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .C1(new_n1036), .C2(new_n1040), .ZN(G57));
endmodule


