//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT21), .B(G898), .Z(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT92), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(G214), .B1(G237), .B2(G902), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G116), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G119), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT5), .ZN(new_n204));
  OAI21_X1  g018(.A(G113), .B1(new_n201), .B2(KEYINPUT5), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n199), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT2), .A2(G113), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT2), .A2(G113), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(KEYINPUT64), .A2(KEYINPUT2), .A3(G113), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT5), .ZN(new_n216));
  OR3_X1    g030(.A1(new_n202), .A2(KEYINPUT5), .A3(G119), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT88), .A4(G113), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n206), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(G104), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT81), .A3(G107), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n221), .A2(G104), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n221), .A2(KEYINPUT3), .A3(G104), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(new_n221), .B2(G104), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n229), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n198), .B1(new_n219), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n227), .A2(new_n233), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n217), .A3(G113), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n237), .A2(new_n199), .B1(new_n214), .B2(new_n208), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n236), .A2(new_n238), .A3(KEYINPUT89), .A4(new_n218), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT80), .A3(G101), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n224), .B2(G107), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n221), .A2(KEYINPUT3), .A3(G104), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n228), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n246), .B2(new_n230), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n246), .B2(new_n230), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n246), .A2(new_n230), .ZN(new_n251));
  INV_X1    g065(.A(new_n213), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n253));
  OAI22_X1  g067(.A1(new_n252), .A2(new_n253), .B1(KEYINPUT2), .B2(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n207), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n248), .A2(new_n251), .B1(new_n255), .B2(new_n215), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n235), .A2(new_n239), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G110), .B(G122), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n197), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n235), .A2(new_n239), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n250), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n258), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  INV_X1    g081(.A(G146), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G143), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT0), .ZN(new_n270));
  INV_X1    g084(.A(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  OAI22_X1  g087(.A1(new_n267), .A2(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n266), .A2(G146), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n275), .B(new_n276), .C1(new_n270), .C2(new_n271), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G125), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G128), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n271), .A2(new_n267), .B1(new_n269), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n275), .A3(new_n276), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G125), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n188), .A2(G224), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n262), .A2(new_n197), .A3(new_n263), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n265), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n215), .A2(new_n237), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n236), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n258), .B(KEYINPUT8), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n295), .B(new_n296), .C1(new_n236), .C2(new_n219), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n279), .A2(new_n287), .A3(new_n298), .A4(new_n289), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n289), .A2(new_n298), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n290), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n257), .A2(new_n258), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n292), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n293), .B1(new_n292), .B2(new_n304), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n195), .B(new_n196), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n308));
  AOI21_X1  g122(.A(G140), .B1(KEYINPUT72), .B2(G125), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n310), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G146), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT72), .A2(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n312), .ZN(new_n318));
  NAND3_X1  g132(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(KEYINPUT16), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n268), .A3(new_n314), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(G237), .ZN(new_n325));
  INV_X1    g139(.A(G237), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT66), .ZN(new_n327));
  OAI211_X1 g141(.A(G214), .B(new_n188), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n266), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(KEYINPUT66), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(G237), .ZN(new_n331));
  AOI21_X1  g145(.A(G953), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G143), .A3(G214), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n323), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n322), .B1(new_n334), .B2(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  AND4_X1   g150(.A1(G143), .A2(new_n336), .A3(G214), .A4(new_n188), .ZN(new_n337));
  AOI21_X1  g151(.A(G143), .B1(new_n332), .B2(G214), .ZN(new_n338));
  OAI21_X1  g152(.A(G131), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n329), .A2(new_n323), .A3(new_n333), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n224), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT18), .B(G131), .C1(new_n337), .C2(new_n338), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n318), .A2(G146), .A3(new_n319), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n286), .A2(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n313), .A2(new_n348), .A3(new_n268), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT18), .A2(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n329), .A2(new_n333), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n343), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n352), .A2(new_n350), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n339), .A2(new_n341), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n268), .B1(new_n320), .B2(new_n314), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n318), .A2(KEYINPUT19), .A3(new_n319), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT19), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n313), .A2(new_n348), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT90), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n318), .A2(new_n362), .A3(KEYINPUT19), .A4(new_n319), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n364), .B2(new_n268), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n346), .A2(new_n355), .B1(new_n356), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n345), .B1(new_n366), .B2(KEYINPUT91), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n337), .A2(new_n338), .A3(G131), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n365), .B1(new_n368), .B2(new_n334), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT91), .B1(new_n369), .B2(new_n353), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n354), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G475), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n343), .A2(new_n345), .A3(new_n353), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(KEYINPUT91), .A3(new_n353), .ZN(new_n377));
  INV_X1    g191(.A(new_n345), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n379), .B2(new_n370), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n373), .ZN(new_n382));
  INV_X1    g196(.A(G902), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n345), .B1(new_n343), .B2(new_n353), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n354), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n375), .A2(new_n382), .B1(G475), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n266), .A2(G128), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n271), .A2(G143), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G134), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G116), .B(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n221), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n202), .A2(KEYINPUT14), .A3(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n392), .ZN(new_n395));
  OAI211_X1 g209(.A(G107), .B(new_n394), .C1(new_n395), .C2(KEYINPUT14), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n387), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n388), .B1(new_n398), .B2(KEYINPUT13), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G134), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n392), .B(new_n221), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n389), .A2(new_n390), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT9), .B(G234), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(G953), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n397), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n397), .B2(new_n405), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n383), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G478), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(KEYINPUT15), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n411), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n386), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n307), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G221), .B1(new_n406), .B2(G902), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n251), .A2(new_n248), .B1(new_n274), .B2(new_n277), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n250), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n284), .A2(KEYINPUT82), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n283), .A2(new_n275), .A3(new_n276), .A4(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n422), .A2(new_n282), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n421), .B1(new_n425), .B2(new_n234), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n285), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n390), .B2(G137), .ZN(new_n430));
  INV_X1    g244(.A(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT11), .A3(G134), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n390), .A2(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n432), .A3(new_n323), .A4(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT83), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  INV_X1    g254(.A(G227), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n428), .A2(KEYINPUT84), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n420), .A2(new_n426), .A3(new_n448), .A4(new_n427), .ZN(new_n449));
  AND4_X1   g263(.A1(new_n446), .A2(new_n447), .A3(new_n437), .A4(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n437), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n428), .B2(KEYINPUT84), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n446), .B1(new_n452), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n445), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n234), .A2(new_n284), .A3(new_n282), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n234), .B2(new_n425), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n437), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(KEYINPUT12), .A3(new_n437), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n444), .B1(new_n461), .B2(new_n439), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n454), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G469), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT86), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT86), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n447), .A2(new_n437), .A3(new_n449), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT85), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n452), .A2(new_n446), .A3(new_n449), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n462), .B1(new_n471), .B2(new_n445), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n467), .B(G469), .C1(new_n472), .C2(G902), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT87), .B(G469), .Z(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n444), .B1(new_n471), .B2(new_n439), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n461), .A2(new_n439), .A3(new_n444), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n383), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n466), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n417), .A2(new_n418), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n407), .B1(G234), .B2(new_n383), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n200), .B2(G128), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT23), .ZN(new_n485));
  INV_X1    g299(.A(G110), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n200), .A2(G128), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n483), .B(new_n488), .C1(new_n200), .C2(G128), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n271), .A2(G119), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT69), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n493), .A2(new_n487), .A3(KEYINPUT69), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n486), .A2(KEYINPUT24), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G110), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT70), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT70), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  OAI22_X1  g314(.A1(new_n494), .A2(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n484), .A2(KEYINPUT23), .B1(new_n200), .B2(G128), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(KEYINPUT73), .A3(new_n486), .A4(new_n489), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n316), .A2(new_n349), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n495), .A2(new_n494), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(G110), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n322), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT74), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n504), .A2(new_n505), .B1(new_n510), .B2(new_n322), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n506), .A2(new_n511), .A3(new_n515), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT75), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n524), .A3(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n526), .A3(new_n383), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT25), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n520), .A2(new_n517), .B1(new_n523), .B2(new_n525), .ZN(new_n531));
  INV_X1    g345(.A(new_n529), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n383), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n482), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n531), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n481), .A2(G902), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT77), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT78), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n531), .B2(new_n383), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n383), .A2(new_n521), .A3(new_n526), .A4(new_n532), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n481), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n543));
  INV_X1    g357(.A(new_n538), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n390), .A2(G137), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n431), .A2(G134), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n283), .A2(new_n275), .A3(new_n276), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n271), .A2(new_n268), .A3(G143), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n283), .B2(new_n276), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n436), .B(new_n550), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n435), .A2(new_n436), .B1(new_n274), .B2(new_n277), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n547), .B(KEYINPUT30), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n437), .A2(new_n278), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n547), .A2(KEYINPUT30), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n547), .A2(KEYINPUT30), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n558), .A2(new_n559), .A3(new_n554), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n255), .A2(new_n215), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n255), .A2(new_n215), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n558), .A2(new_n566), .A3(new_n554), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n332), .A2(G210), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT27), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT26), .B(G101), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n564), .A2(new_n565), .A3(new_n567), .A4(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT67), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n567), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n562), .B2(new_n563), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(KEYINPUT67), .A3(new_n565), .A4(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n570), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n569), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT28), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n563), .B1(new_n555), .B2(new_n556), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n567), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n555), .A2(new_n556), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT28), .B1(new_n584), .B2(new_n566), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n580), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n565), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n576), .A2(new_n571), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G472), .A2(G902), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT68), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT68), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n574), .A2(new_n577), .B1(new_n588), .B2(new_n587), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT32), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G472), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n580), .A2(new_n583), .A3(new_n585), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(KEYINPUT29), .ZN(new_n601));
  INV_X1    g415(.A(new_n576), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n580), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n600), .B2(KEYINPUT29), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n594), .A2(new_n595), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(KEYINPUT32), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n546), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n546), .A2(new_n609), .A3(KEYINPUT79), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n480), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n230), .ZN(G3));
  NAND2_X1  g429(.A1(new_n479), .A2(new_n418), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT68), .B1(new_n590), .B2(new_n591), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n594), .A2(new_n593), .A3(new_n595), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n594), .B2(G902), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n539), .A3(new_n545), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n385), .A2(G475), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n380), .A2(new_n381), .A3(new_n373), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n381), .B1(new_n380), .B2(new_n373), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OR3_X1    g440(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT33), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT33), .B1(new_n409), .B2(new_n410), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(G478), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(G478), .A2(G902), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n629), .B(new_n630), .C1(G478), .C2(new_n411), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT93), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT93), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n635), .A3(new_n632), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n307), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AOI21_X1  g454(.A(new_n415), .B1(new_n375), .B2(new_n382), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n316), .A2(new_n321), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n339), .B2(new_n340), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n353), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n378), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n646), .B2(new_n376), .ZN(new_n647));
  INV_X1    g461(.A(G475), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(KEYINPUT94), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT94), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n385), .B2(G475), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n641), .A2(KEYINPUT95), .A3(new_n652), .A4(new_n195), .ZN(new_n653));
  INV_X1    g467(.A(new_n196), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n292), .A2(new_n304), .ZN(new_n655));
  INV_X1    g469(.A(new_n293), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n292), .A2(new_n293), .A3(new_n304), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n414), .B1(new_n624), .B2(new_n625), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT94), .B1(new_n647), .B2(new_n648), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n385), .A2(new_n650), .A3(G475), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT95), .B1(new_n665), .B2(new_n195), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n622), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  AND2_X1   g484(.A1(new_n479), .A2(new_n418), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n592), .A2(new_n596), .A3(new_n620), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n512), .B(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n537), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n542), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n671), .A2(new_n417), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT96), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT37), .B(G110), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  XOR2_X1   g497(.A(new_n189), .B(KEYINPUT97), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(new_n193), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n659), .A2(new_n665), .A3(KEYINPUT98), .A4(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT98), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n375), .A2(new_n382), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n652), .A2(new_n691), .A3(new_n414), .A4(new_n688), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n196), .B1(new_n305), .B2(new_n306), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n609), .A2(new_n479), .A3(new_n418), .A4(new_n677), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT99), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n609), .A2(new_n479), .A3(new_n418), .A4(new_n677), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT99), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n689), .A2(new_n694), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n602), .A2(new_n571), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n582), .A2(new_n567), .ZN(new_n706));
  AOI21_X1  g520(.A(G902), .B1(new_n580), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n599), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n607), .B2(KEYINPUT32), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n598), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n704), .B1(new_n598), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n657), .A2(new_n658), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n415), .A2(new_n654), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n626), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n678), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n687), .B(KEYINPUT39), .Z(new_n718));
  AND2_X1   g532(.A1(new_n671), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n719), .A2(KEYINPUT40), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(KEYINPUT40), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n712), .B(new_n717), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n266), .ZN(G45));
  NAND3_X1  g537(.A1(new_n626), .A2(new_n632), .A3(new_n688), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT101), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n626), .A2(new_n726), .A3(new_n632), .A4(new_n688), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n659), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(KEYINPUT102), .A3(new_n659), .A4(new_n727), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n698), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NAND2_X1  g547(.A1(new_n539), .A2(new_n545), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n598), .B2(new_n608), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n439), .B1(new_n450), .B2(new_n453), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n477), .B1(new_n736), .B2(new_n443), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(G902), .A3(new_n474), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n443), .ZN(new_n739));
  INV_X1    g553(.A(new_n477), .ZN(new_n740));
  AOI21_X1  g554(.A(G902), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n465), .B1(new_n741), .B2(KEYINPUT103), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n737), .B2(G902), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n738), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n735), .A2(new_n418), .A3(new_n745), .A4(new_n637), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  OAI211_X1 g562(.A(KEYINPUT103), .B(new_n383), .C1(new_n476), .C2(new_n477), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n744), .A2(new_n749), .A3(G469), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n750), .A2(new_n418), .A3(new_n478), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n667), .A3(new_n735), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  AND4_X1   g567(.A1(new_n418), .A2(new_n750), .A3(new_n478), .A4(new_n659), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n416), .A2(new_n194), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n609), .A2(new_n755), .A3(new_n677), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G119), .ZN(G21));
  INV_X1    g572(.A(KEYINPUT104), .ZN(new_n759));
  AOI21_X1  g573(.A(G902), .B1(new_n578), .B2(new_n589), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n759), .B1(new_n760), .B2(new_n599), .ZN(new_n761));
  INV_X1    g575(.A(new_n607), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n542), .A2(new_n544), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT104), .B(G472), .C1(new_n594), .C2(G902), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n716), .A2(new_n195), .A3(new_n713), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n751), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  NAND4_X1  g584(.A1(new_n761), .A2(new_n677), .A3(new_n762), .A4(new_n765), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n725), .A2(KEYINPUT105), .A3(new_n727), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n631), .B1(new_n691), .B2(new_n623), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n726), .B1(new_n775), .B2(new_n688), .ZN(new_n776));
  INV_X1    g590(.A(new_n727), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n754), .A2(new_n772), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n418), .A2(new_n196), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n305), .A2(new_n306), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n464), .A2(new_n465), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(new_n738), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n778), .A2(new_n735), .A3(new_n773), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n725), .A2(KEYINPUT105), .A3(new_n727), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT105), .B1(new_n725), .B2(new_n727), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n610), .A2(new_n786), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT106), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n781), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n788), .A2(new_n789), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(KEYINPUT106), .A3(new_n794), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT107), .A4(new_n782), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n762), .A2(new_n597), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n764), .B1(new_n801), .B2(new_n608), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n793), .A2(KEYINPUT42), .A3(new_n787), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  XNOR2_X1  g619(.A(new_n692), .B(KEYINPUT108), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n735), .A2(new_n806), .A3(new_n787), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G134), .ZN(G36));
  NAND3_X1  g622(.A1(new_n657), .A2(new_n196), .A3(new_n658), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT109), .Z(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n386), .A2(new_n632), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(new_n672), .A3(new_n677), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n811), .B1(new_n815), .B2(KEYINPUT44), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT110), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n672), .A3(new_n677), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(KEYINPUT110), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n472), .A2(KEYINPUT45), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n472), .A2(KEYINPUT45), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(G469), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(G469), .A2(G902), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n738), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n829), .A2(new_n418), .A3(new_n718), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n817), .A2(new_n820), .A3(new_n821), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  INV_X1    g646(.A(new_n809), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n725), .A2(new_n734), .A3(new_n727), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n609), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n829), .A2(KEYINPUT47), .A3(new_n418), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT47), .B1(new_n829), .B2(new_n418), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  OAI211_X1 g653(.A(new_n623), .B(new_n414), .C1(new_n624), .C2(new_n625), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n691), .A2(new_n842), .A3(new_n623), .A4(new_n414), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n307), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT111), .B1(new_n307), .B2(new_n633), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n659), .A2(new_n775), .A3(new_n848), .A4(new_n195), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n622), .A2(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n752), .A2(new_n851), .A3(new_n757), .A4(new_n769), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n786), .A2(new_n771), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n778), .A2(new_n853), .A3(new_n773), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n678), .B1(new_n598), .B2(new_n608), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n691), .A2(new_n415), .A3(new_n688), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n809), .A2(new_n856), .A3(new_n664), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n671), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n807), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n746), .A2(new_n680), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n614), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n854), .A2(new_n807), .A3(new_n858), .A4(KEYINPUT113), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n852), .A2(new_n861), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n800), .B2(new_n803), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT99), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n779), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n713), .A2(new_n626), .A3(new_n715), .ZN(new_n871));
  INV_X1    g685(.A(new_n418), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n677), .A2(new_n872), .A3(new_n687), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n478), .B1(new_n465), .B2(new_n464), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n710), .B2(new_n711), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n732), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n869), .A2(new_n870), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n791), .A2(new_n792), .A3(new_n771), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n701), .A2(new_n697), .B1(new_n879), .B2(new_n754), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n732), .A2(new_n876), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT52), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT116), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n870), .B1(new_n869), .B2(new_n877), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n881), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n866), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n869), .B2(new_n877), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT115), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n892), .C1(new_n869), .C2(new_n877), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n896), .A3(new_n886), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT53), .B1(new_n897), .B2(new_n866), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n888), .A2(new_n889), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(KEYINPUT53), .A3(new_n866), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n814), .A2(new_n767), .A3(new_n685), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n714), .A2(new_n196), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n751), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT50), .Z(new_n908));
  AND2_X1   g722(.A1(new_n751), .A2(new_n833), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n712), .A3(new_n546), .A4(new_n189), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n910), .A2(new_n626), .A3(new_n632), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n909), .A2(new_n685), .A3(new_n814), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n772), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n908), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n836), .A2(new_n837), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n745), .A2(new_n872), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n905), .A2(new_n810), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT51), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT51), .A4(new_n913), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n915), .A2(KEYINPUT117), .A3(new_n916), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n922), .A2(new_n918), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n912), .A2(new_n802), .ZN(new_n927));
  XOR2_X1   g741(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n188), .A2(G952), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n905), .B2(new_n754), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n634), .A2(new_n636), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n929), .B(new_n931), .C1(new_n933), .C2(new_n910), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n920), .A2(new_n926), .A3(new_n934), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n904), .A2(new_n935), .B1(G952), .B2(G953), .ZN(new_n936));
  INV_X1    g750(.A(new_n745), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT49), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT49), .ZN(new_n939));
  NOR4_X1   g753(.A1(new_n714), .A2(new_n764), .A3(new_n783), .A4(new_n812), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n938), .A2(new_n712), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n936), .A2(new_n941), .ZN(G75));
  NAND2_X1  g756(.A1(new_n265), .A2(new_n291), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n290), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT55), .Z(new_n945));
  INV_X1    g759(.A(G210), .ZN(new_n946));
  AOI211_X1 g760(.A(new_n946), .B(new_n383), .C1(new_n900), .C2(new_n902), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n947), .B2(KEYINPUT56), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  INV_X1    g763(.A(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n900), .A2(new_n902), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(G902), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n949), .B(new_n950), .C1(new_n952), .C2(new_n946), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n188), .A2(G952), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n948), .A2(new_n953), .A3(new_n955), .ZN(G51));
  XOR2_X1   g770(.A(new_n825), .B(KEYINPUT57), .Z(new_n957));
  AND3_X1   g771(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n737), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n952), .A2(new_n824), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(G54));
  NAND2_X1  g778(.A1(KEYINPUT58), .A2(G475), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n383), .B(new_n965), .C1(new_n900), .C2(new_n902), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT119), .B1(new_n966), .B2(new_n380), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n954), .B1(new_n966), .B2(new_n380), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n969), .B(new_n372), .C1(new_n952), .C2(new_n965), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(new_n627), .A2(new_n628), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT120), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n630), .B(KEYINPUT59), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n974), .C1(new_n958), .C2(new_n959), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n955), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n904), .B2(new_n974), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G63));
  XNOR2_X1  g792(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n900), .B2(new_n902), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n674), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n531), .B(KEYINPUT122), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n955), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n979), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n900), .A2(new_n902), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n989), .B2(new_n981), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(KEYINPUT61), .A3(new_n955), .A4(new_n983), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(G66));
  INV_X1    g806(.A(G224), .ZN(new_n993));
  OAI21_X1  g807(.A(G953), .B1(new_n192), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n852), .A2(new_n863), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n943), .B1(G898), .B2(new_n188), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT123), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(G69));
  XOR2_X1   g814(.A(new_n364), .B(KEYINPUT124), .Z(new_n1001));
  XNOR2_X1  g815(.A(new_n562), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G900), .A2(G953), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n802), .A2(new_n871), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n830), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n831), .A2(new_n807), .A3(new_n838), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n804), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n880), .A2(new_n732), .ZN(new_n1008));
  OR3_X1    g822(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1002), .B(new_n1003), .C1(new_n1009), .C2(G953), .ZN(new_n1010));
  OAI21_X1  g824(.A(G953), .B1(new_n441), .B2(new_n686), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n1002), .B2(KEYINPUT126), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n612), .A2(new_n613), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n841), .A2(new_n843), .A3(new_n633), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1014), .A2(new_n719), .A3(new_n833), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n830), .B1(KEYINPUT110), .B2(new_n816), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n821), .A2(new_n820), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(KEYINPUT125), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT125), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n831), .A2(new_n1021), .A3(new_n1016), .ZN(new_n1022));
  INV_X1    g836(.A(new_n915), .ZN(new_n1023));
  AOI22_X1  g837(.A1(new_n1020), .A2(new_n1022), .B1(new_n1023), .B2(new_n835), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n722), .A2(new_n1008), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1028), .A2(new_n188), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1010), .B(new_n1013), .C1(new_n1029), .C2(new_n1002), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1010), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1002), .B1(new_n1028), .B2(new_n188), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1012), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1030), .A2(new_n1033), .ZN(G72));
  NAND4_X1  g848(.A1(new_n1024), .A2(new_n1026), .A3(new_n996), .A4(new_n1027), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  NAND2_X1  g851(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n705), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n954), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n602), .A2(new_n571), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1037), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1043), .B1(new_n890), .B2(new_n898), .ZN(new_n1044));
  OAI211_X1 g858(.A(KEYINPUT127), .B(new_n1037), .C1(new_n1009), .C2(new_n995), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT127), .ZN(new_n1046));
  NOR4_X1   g860(.A1(new_n1006), .A2(new_n1007), .A3(new_n995), .A4(new_n1008), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1046), .B1(new_n1047), .B2(new_n1042), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1045), .A2(new_n1048), .A3(new_n1041), .ZN(new_n1049));
  AND3_X1   g863(.A1(new_n1040), .A2(new_n1044), .A3(new_n1049), .ZN(G57));
endmodule


