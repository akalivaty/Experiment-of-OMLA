//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n209), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G87), .A2(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n205), .C2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n225), .B(new_n230), .C1(G50), .C2(G226), .ZN(new_n231));
  AND2_X1   g0031(.A1(KEYINPUT65), .A2(G77), .ZN(new_n232));
  NOR2_X1   g0032(.A1(KEYINPUT65), .A2(G77), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G244), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n221), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(KEYINPUT1), .ZN(new_n238));
  OAI21_X1  g0038(.A(new_n220), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n213), .B(new_n239), .C1(new_n238), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n228), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT66), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT8), .B(G58), .Z(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n218), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT15), .B(G87), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n260), .B1(new_n218), .B2(new_n234), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n217), .B1(new_n209), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(new_n267), .A3(G13), .A4(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n265), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G77), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n271), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n234), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n266), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n264), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n279), .ZN(new_n285));
  INV_X1    g0085(.A(G244), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(G1698), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n290), .B1(new_n206), .B2(new_n288), .C1(new_n291), .C2(new_n224), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G169), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n257), .B1(new_n278), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n266), .A2(new_n274), .A3(new_n277), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(KEYINPUT70), .C1(G169), .C2(new_n294), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n294), .A2(G190), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n278), .B(new_n302), .C1(new_n303), .C2(new_n294), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n289), .A2(G222), .ZN(new_n306));
  AND2_X1   g0106(.A1(G223), .A2(G1698), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n288), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n234), .B2(new_n288), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT67), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n284), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n310), .B2(new_n309), .ZN(new_n312));
  INV_X1    g0112(.A(new_n285), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n281), .B1(new_n313), .B2(G226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n299), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n272), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n272), .A2(new_n318), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n273), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n202), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(new_n261), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n265), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(G50), .B2(new_n275), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n315), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n317), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n316), .A2(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(KEYINPUT9), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n315), .B2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT9), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n322), .B2(new_n328), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n305), .B(new_n333), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n276), .A2(new_n223), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  INV_X1    g0145(.A(new_n259), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n202), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n261), .A2(new_n348), .B1(new_n218), .B2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n265), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT11), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n272), .A2(G68), .A3(new_n273), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n288), .A2(new_n289), .ZN(new_n356));
  INV_X1    g0156(.A(G226), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n293), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n281), .B1(new_n313), .B2(G238), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT13), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(KEYINPUT14), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT14), .B1(new_n365), .B2(new_n366), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n365), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT73), .B1(new_n365), .B2(new_n299), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n353), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n365), .A2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(new_n353), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(new_n365), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n357), .A2(G1698), .ZN(new_n380));
  AND2_X1   g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n380), .B1(G223), .B2(G1698), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT75), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n284), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n384), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n282), .B1(new_n285), .B2(new_n228), .ZN(new_n389));
  OAI21_X1  g0189(.A(G200), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G190), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(G58), .B(G68), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n381), .A2(new_n382), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n288), .B2(G20), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT74), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n218), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n399), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n398), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT16), .B(new_n395), .C1(new_n405), .C2(new_n223), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n400), .A2(new_n397), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n395), .B1(new_n407), .B2(new_n223), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n410), .A3(new_n265), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n321), .A2(new_n258), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n275), .A2(new_n323), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n393), .A2(KEYINPUT17), .A3(new_n411), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n414), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n391), .A2(G179), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n331), .B2(new_n391), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n421), .A3(new_n418), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n411), .A2(new_n390), .A3(new_n414), .A4(new_n392), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n415), .A2(new_n420), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n343), .A2(new_n379), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G87), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n429), .A2(KEYINPUT81), .A3(G20), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n288), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT22), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n218), .A2(G107), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT23), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G116), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n434), .A2(new_n435), .B1(G20), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n288), .A2(KEYINPUT22), .A3(new_n430), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n434), .A2(new_n440), .A3(new_n435), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n435), .A2(new_n206), .A3(G20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n433), .A2(new_n438), .A3(new_n439), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT24), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n444), .A2(new_n439), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT24), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n437), .B1(new_n431), .B2(new_n432), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n327), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n276), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT25), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n275), .B2(G107), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n264), .A2(G1), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT76), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n272), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(new_n206), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n267), .A2(G45), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(KEYINPUT77), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT77), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n466));
  AOI21_X1  g0266(.A(G41), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g0269(.A(KEYINPUT78), .B(G41), .C1(new_n464), .C2(new_n466), .ZN(new_n470));
  OAI211_X1 g0270(.A(G264), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n288), .A2(G250), .A3(new_n289), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n288), .A2(G257), .A3(G1698), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n293), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n464), .A2(new_n466), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT78), .B1(new_n477), .B2(G41), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n467), .A2(new_n468), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n293), .A2(new_n280), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n463), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n471), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G200), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n460), .B(new_n483), .C1(new_n377), .C2(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n331), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n471), .A2(new_n476), .A3(new_n481), .A4(new_n299), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n451), .C2(new_n459), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n445), .A2(KEYINPUT24), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n265), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n458), .A2(new_n206), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n454), .B2(new_n452), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(new_n486), .A4(new_n485), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(new_n488), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n498), .A2(new_n205), .A3(G107), .ZN(new_n499));
  XNOR2_X1  g0299(.A(G97), .B(G107), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(new_n218), .B1(new_n348), .B2(new_n346), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n206), .B1(new_n400), .B2(new_n397), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n265), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n457), .A2(new_n272), .A3(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n276), .A2(new_n205), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G244), .B(new_n289), .C1(new_n381), .C2(new_n382), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n289), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n293), .ZN(new_n516));
  OAI211_X1 g0316(.A(G257), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n481), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n508), .B1(G200), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n518), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n518), .A2(new_n331), .B1(new_n504), .B2(new_n507), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n516), .A2(new_n299), .A3(new_n517), .A4(new_n481), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n218), .B1(new_n355), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G87), .B2(new_n207), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n261), .B2(new_n205), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n218), .B(G68), .C1(new_n381), .C2(new_n382), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n265), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n276), .A2(new_n262), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n457), .A2(new_n272), .A3(G87), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n461), .A2(G250), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n293), .A2(new_n537), .B1(new_n280), .B2(new_n461), .ZN(new_n538));
  OAI211_X1 g0338(.A(G238), .B(new_n289), .C1(new_n381), .C2(new_n382), .ZN(new_n539));
  OAI211_X1 g0339(.A(G244), .B(G1698), .C1(new_n381), .C2(new_n382), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n436), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n293), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(G190), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n531), .A2(new_n265), .B1(new_n276), .B2(new_n262), .ZN(new_n547));
  INV_X1    g0347(.A(new_n262), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n457), .A2(new_n272), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(new_n549), .B1(new_n542), .B2(new_n299), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n331), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n522), .A2(new_n525), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n497), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT80), .ZN(new_n556));
  OAI211_X1 g0356(.A(G270), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n481), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(KEYINPUT79), .A3(new_n481), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  OAI221_X1 g0364(.A(new_n563), .B1(new_n229), .B2(new_n356), .C1(new_n564), .C2(new_n288), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n293), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n556), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n557), .A2(KEYINPUT79), .A3(new_n481), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT79), .B1(new_n557), .B2(new_n481), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n556), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(G190), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n276), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n458), .B2(new_n573), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n513), .B(new_n218), .C1(G33), .C2(new_n205), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(new_n265), .C1(new_n218), .C2(G116), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT20), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(G200), .A3(new_n570), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n572), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n579), .A2(new_n331), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(KEYINPUT21), .A3(new_n570), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n570), .A3(new_n584), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n562), .A2(G179), .A3(new_n566), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n579), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n586), .A2(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n555), .A2(new_n583), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n428), .A2(new_n592), .ZN(G372));
  INV_X1    g0393(.A(new_n333), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n420), .A2(new_n422), .ZN(new_n595));
  INV_X1    g0395(.A(new_n370), .ZN(new_n596));
  INV_X1    g0396(.A(new_n373), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n301), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n353), .B1(new_n378), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n415), .A2(new_n425), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n341), .A2(new_n342), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n594), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n523), .A2(new_n524), .A3(new_n546), .A4(new_n552), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT26), .ZN(new_n606));
  INV_X1    g0406(.A(new_n538), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n541), .A2(new_n608), .A3(new_n293), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(new_n541), .B2(new_n293), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n331), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n550), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(G200), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n377), .B(new_n538), .C1(new_n293), .C2(new_n541), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n535), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n550), .A2(new_n612), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n518), .A2(new_n331), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n618), .A2(new_n524), .A3(new_n508), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n606), .B(new_n613), .C1(new_n620), .C2(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n586), .A2(new_n587), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n589), .A2(new_n590), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n585), .A3(new_n623), .A4(new_n487), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n484), .A2(new_n525), .A3(new_n522), .A4(new_n617), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n604), .B1(new_n428), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g0427(.A(new_n627), .B(KEYINPUT85), .Z(G369));
  NAND2_X1  g0428(.A1(new_n591), .A2(new_n585), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n267), .A2(new_n218), .A3(G13), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n579), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n629), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n622), .A2(new_n585), .A3(new_n623), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n583), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n640), .B2(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n487), .A2(new_n636), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT86), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n460), .A2(new_n636), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n497), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n635), .B1(new_n591), .B2(new_n585), .ZN(new_n649));
  INV_X1    g0449(.A(new_n487), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n647), .A2(new_n649), .B1(new_n650), .B2(new_n636), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(G399));
  NOR3_X1   g0452(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n210), .A2(new_n283), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(G1), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n215), .B2(new_n654), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT28), .ZN(new_n657));
  INV_X1    g0457(.A(G330), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n520), .A2(new_n471), .A3(new_n476), .A4(new_n542), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT30), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n588), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n588), .B2(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n581), .A2(new_n570), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n518), .A2(new_n611), .A3(new_n299), .A4(new_n482), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n635), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n592), .B2(new_n635), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT31), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT31), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n658), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT29), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT87), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n613), .B1(new_n605), .B2(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n617), .B2(new_n619), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n674), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n614), .A2(new_n616), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n613), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT26), .B1(new_n680), .B2(new_n525), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n553), .A2(new_n619), .A3(new_n676), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n681), .A2(KEYINPUT87), .A3(new_n682), .A4(new_n613), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n488), .A2(new_n496), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n622), .A2(new_n685), .A3(new_n585), .A4(new_n623), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n625), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n673), .B1(new_n688), .B2(new_n636), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n626), .A2(KEYINPUT29), .A3(new_n635), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n672), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n657), .B1(new_n693), .B2(G1), .ZN(G364));
  OR2_X1    g0494(.A1(new_n641), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(G13), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G20), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n267), .B1(new_n697), .B2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n654), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n695), .A2(new_n642), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT88), .ZN(new_n704));
  NOR2_X1   g0504(.A1(G13), .A2(G33), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT89), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT92), .Z(new_n708));
  NOR2_X1   g0508(.A1(new_n641), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n217), .B1(G20), .B2(new_n331), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n288), .A2(new_n210), .ZN(new_n713));
  INV_X1    g0513(.A(G355), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(G116), .B2(new_n210), .ZN(new_n715));
  INV_X1    g0515(.A(G45), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n251), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n396), .A2(new_n210), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n716), .B2(new_n216), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n218), .A2(G190), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G159), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT32), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n303), .A2(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n206), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n396), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n299), .A2(new_n303), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n731), .A2(new_n721), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n218), .A2(new_n377), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n727), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n730), .B1(new_n223), .B2(new_n733), .C1(new_n429), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n722), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n726), .B(new_n736), .C1(G97), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n299), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n721), .A2(new_n740), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(G58), .A2(new_n742), .B1(new_n744), .B2(new_n235), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n731), .A2(new_n734), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n202), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT90), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n741), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  INV_X1    g0552(.A(G329), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n728), .A2(new_n752), .B1(new_n723), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n751), .B(new_n754), .C1(G326), .C2(new_n746), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n735), .A2(new_n564), .B1(new_n743), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  OAI21_X1  g0558(.A(new_n396), .B1(new_n733), .B2(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n757), .B(new_n759), .C1(G294), .C2(new_n738), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n739), .A2(new_n749), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n710), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n701), .B1(new_n712), .B2(new_n720), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT91), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n709), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n704), .A2(new_n765), .ZN(G396));
  NAND2_X1  g0566(.A1(new_n624), .A2(new_n625), .ZN(new_n767));
  INV_X1    g0567(.A(new_n621), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n635), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT95), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n301), .A2(new_n304), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n297), .A2(new_n635), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n301), .A2(new_n770), .A3(new_n297), .A4(new_n635), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(KEYINPUT96), .B1(new_n769), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT96), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n626), .A2(new_n778), .A3(new_n775), .A4(new_n635), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n775), .B1(new_n626), .B2(new_n635), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n701), .B1(new_n782), .B2(new_n672), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n672), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n710), .A2(new_n705), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n702), .B1(new_n348), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G143), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n741), .A2(new_n787), .B1(new_n743), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n733), .A2(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n789), .B(new_n791), .C1(G137), .C2(new_n746), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n288), .B1(new_n728), .B2(new_n223), .ZN(new_n795));
  INV_X1    g0595(.A(G132), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n735), .A2(new_n202), .B1(new_n723), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(G58), .C2(new_n738), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n793), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n728), .A2(new_n429), .B1(new_n723), .B2(new_n756), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n747), .A2(new_n564), .B1(new_n741), .B2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(G97), .C2(new_n738), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n396), .B1(new_n735), .B2(new_n206), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G116), .A2(new_n744), .B1(new_n732), .B2(G283), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n803), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n799), .A2(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n786), .B1(new_n762), .B2(new_n809), .C1(new_n776), .C2(new_n706), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n784), .A2(new_n810), .ZN(G384));
  NOR2_X1   g0611(.A1(new_n697), .A2(new_n267), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n353), .A2(new_n635), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n596), .B2(new_n597), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n374), .A2(new_n378), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n639), .A2(new_n583), .A3(new_n555), .A4(new_n636), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n669), .B1(new_n818), .B2(new_n666), .ZN(new_n819));
  INV_X1    g0619(.A(new_n670), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n817), .B(new_n776), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n419), .A2(new_n423), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT98), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT37), .ZN(new_n824));
  INV_X1    g0624(.A(new_n633), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n416), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n419), .A2(new_n826), .A3(new_n824), .A4(new_n423), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT98), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n419), .A2(new_n826), .A3(new_n423), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT37), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n827), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n426), .A2(new_n416), .A3(new_n825), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n406), .A2(new_n265), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n395), .B1(new_n405), .B2(new_n223), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n409), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n837), .A2(new_n839), .B1(new_n412), .B2(new_n413), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n423), .B1(new_n840), .B2(new_n633), .ZN(new_n841));
  OAI21_X1  g0641(.A(G169), .B1(new_n388), .B2(new_n389), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n842), .A2(new_n417), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n828), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n840), .A2(new_n633), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n426), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n836), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT40), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT99), .B1(new_n821), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT40), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n846), .A2(new_n848), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n835), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n849), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n853), .B1(new_n821), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n775), .B1(new_n668), .B2(new_n670), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n836), .B2(new_n849), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT99), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n817), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n852), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n427), .B1(new_n819), .B2(new_n820), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n865), .A2(new_n866), .A3(new_n658), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n832), .B2(new_n833), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n374), .A2(new_n635), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n849), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n595), .A2(new_n825), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n599), .A2(new_n636), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT97), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n777), .B2(new_n779), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n856), .A3(new_n817), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n427), .B1(new_n689), .B2(new_n690), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n604), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n882), .B(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n812), .B1(new_n868), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n868), .ZN(new_n887));
  INV_X1    g0687(.A(new_n501), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(KEYINPUT35), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(KEYINPUT35), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(G116), .A3(new_n219), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n216), .B1(new_n227), .B2(new_n223), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n893), .A2(new_n234), .B1(G50), .B2(new_n223), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n696), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n887), .A2(new_n892), .A3(new_n895), .ZN(G367));
  OAI21_X1  g0696(.A(new_n711), .B1(new_n210), .B2(new_n262), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n247), .A2(new_n718), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n701), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n396), .B1(new_n741), .B2(new_n564), .ZN(new_n900));
  INV_X1    g0700(.A(G317), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n747), .A2(new_n756), .B1(new_n723), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n900), .B(new_n902), .C1(G107), .C2(new_n738), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G283), .A2(new_n744), .B1(new_n732), .B2(G294), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n205), .B2(new_n728), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT102), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n735), .B2(new_n573), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(KEYINPUT46), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n903), .B(new_n908), .C1(KEYINPUT46), .C2(new_n907), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n747), .A2(new_n787), .B1(new_n741), .B2(new_n790), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n733), .A2(new_n788), .B1(new_n234), .B2(new_n728), .ZN(new_n911));
  INV_X1    g0711(.A(new_n738), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n223), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n288), .B1(new_n743), .B2(new_n202), .ZN(new_n914));
  OR4_X1    g0714(.A1(new_n910), .A2(new_n911), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(KEYINPUT103), .B(G137), .Z(new_n916));
  OAI22_X1  g0716(.A1(new_n916), .A2(new_n723), .B1(new_n735), .B2(new_n227), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT104), .Z(new_n918));
  OAI21_X1  g0718(.A(new_n909), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT47), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n899), .B1(new_n920), .B2(new_n710), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n612), .A2(new_n550), .A3(new_n535), .A4(new_n635), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n536), .A2(new_n636), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n680), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(new_n708), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT101), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n647), .A2(new_n649), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n650), .A2(new_n636), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n508), .A2(new_n635), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n522), .A2(new_n525), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n619), .A2(new_n635), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n928), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n651), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(KEYINPUT44), .A3(new_n936), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT44), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n651), .B2(new_n935), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n648), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n648), .B1(new_n939), .B2(new_n943), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n647), .B(new_n649), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n642), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n692), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n654), .B(KEYINPUT41), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n927), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n939), .A2(new_n943), .ZN(new_n954));
  INV_X1    g0754(.A(new_n648), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n956), .A2(new_n693), .A3(new_n944), .A4(new_n950), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n693), .ZN(new_n958));
  INV_X1    g0758(.A(new_n952), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(KEYINPUT101), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n699), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT100), .B(KEYINPUT43), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n924), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT43), .B2(new_n924), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n647), .A2(new_n649), .A3(new_n935), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n525), .B1(new_n685), .B2(new_n933), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n636), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  MUX2_X1   g0770(.A(new_n963), .B(new_n964), .S(new_n970), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n648), .A2(new_n936), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n926), .B1(new_n961), .B2(new_n974), .ZN(G387));
  NAND2_X1  g0775(.A1(new_n693), .A2(new_n950), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n692), .A2(new_n949), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n700), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n647), .A2(new_n708), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n713), .A2(new_n653), .B1(G107), .B2(new_n210), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n244), .A2(new_n716), .ZN(new_n981));
  INV_X1    g0781(.A(new_n653), .ZN(new_n982));
  AOI211_X1 g0782(.A(G45), .B(new_n982), .C1(G68), .C2(G77), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n323), .A2(G50), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT50), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n718), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n980), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n735), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n235), .A2(new_n988), .B1(new_n746), .B2(G159), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n288), .C1(new_n205), .C2(new_n728), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n743), .A2(new_n223), .B1(new_n723), .B2(new_n790), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n733), .A2(new_n323), .B1(new_n202), .B2(new_n741), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n912), .A2(new_n262), .ZN(new_n993));
  NOR4_X1   g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n988), .A2(G294), .B1(new_n738), .B2(G283), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G322), .A2(new_n746), .B1(new_n732), .B2(G311), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n564), .B2(new_n743), .C1(new_n901), .C2(new_n741), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT48), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n998), .B2(new_n997), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT49), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n288), .B1(new_n724), .B2(G326), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n573), .B2(new_n728), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1000), .B2(KEYINPUT49), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n994), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n701), .B1(new_n712), .B2(new_n987), .C1(new_n1005), .C2(new_n762), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT105), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n950), .A2(new_n699), .B1(new_n979), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n978), .A2(new_n1008), .ZN(G393));
  OAI21_X1  g0809(.A(new_n976), .B1(new_n945), .B2(new_n946), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(new_n700), .A3(new_n957), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n936), .A2(new_n707), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n255), .A2(new_n210), .A3(new_n396), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n711), .B1(new_n205), .B2(new_n210), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n701), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n742), .A2(G311), .B1(new_n746), .B2(G317), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT52), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n735), .A2(new_n752), .B1(new_n723), .B2(new_n750), .ZN(new_n1018));
  OR4_X1    g0818(.A1(new_n288), .A2(new_n1017), .A3(new_n729), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n733), .A2(new_n564), .B1(new_n743), .B2(new_n801), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G116), .B2(new_n738), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT108), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G68), .A2(new_n988), .B1(new_n724), .B2(G143), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n288), .C1(new_n429), .C2(new_n728), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT106), .Z(new_n1025));
  OAI22_X1  g0825(.A1(new_n747), .A2(new_n790), .B1(new_n741), .B2(new_n788), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n733), .A2(new_n202), .B1(new_n743), .B2(new_n323), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT107), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(G77), .B2(new_n738), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1027), .B(new_n1030), .C1(new_n1029), .C2(new_n1028), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1019), .A2(new_n1022), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1015), .B1(new_n1032), .B2(new_n710), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n947), .A2(new_n699), .B1(new_n1012), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1011), .A2(new_n1034), .ZN(G390));
  INV_X1    g0835(.A(new_n879), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n635), .B1(new_n684), .B2(new_n687), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n776), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n850), .B1(new_n374), .B2(new_n635), .C1(new_n1038), .C2(new_n816), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n873), .B1(new_n880), .B2(new_n817), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n872), .A2(new_n874), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(G330), .B(new_n776), .C1(new_n819), .C2(new_n820), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n816), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n859), .A2(G330), .A3(new_n817), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n699), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n785), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n701), .B1(new_n258), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n735), .A2(new_n790), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT53), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT54), .B(G143), .ZN(new_n1054));
  INV_X1    g0854(.A(G125), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n743), .A2(new_n1054), .B1(new_n723), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G159), .B2(new_n738), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n288), .B1(new_n728), .B2(new_n202), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT112), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n733), .A2(new_n916), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(KEYINPUT112), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n742), .A2(G132), .B1(new_n746), .B2(G128), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n396), .B1(new_n735), .B2(new_n429), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT113), .Z(new_n1066));
  INV_X1    g0866(.A(new_n728), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G116), .A2(new_n742), .B1(new_n1067), .B2(G68), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G283), .A2(new_n746), .B1(new_n732), .B2(G107), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G97), .A2(new_n744), .B1(new_n724), .B2(G294), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n738), .A2(G77), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1058), .A2(new_n1064), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1051), .B1(new_n1073), .B2(new_n710), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1041), .B2(new_n706), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1048), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(G330), .B(new_n427), .C1(new_n819), .C2(new_n820), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n883), .A2(new_n604), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT109), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n883), .A2(new_n1077), .A3(KEYINPUT109), .A4(new_n604), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n817), .B1(new_n859), .B2(G330), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n880), .B1(new_n1083), .B2(new_n1044), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1043), .A2(new_n816), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1046), .A2(new_n1038), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1045), .A2(new_n1047), .A3(new_n1082), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT110), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1092), .A2(KEYINPUT110), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n654), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1076), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(G378));
  NAND4_X1  g0899(.A1(new_n852), .A2(new_n858), .A3(G330), .A4(new_n862), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n329), .A2(new_n633), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n603), .A2(new_n333), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n603), .B2(new_n333), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(KEYINPUT116), .A3(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n877), .A2(new_n881), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n877), .B2(new_n881), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1101), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1110), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n882), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n877), .A2(new_n881), .A3(new_n1110), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1100), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n706), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1108), .A2(new_n1123), .A3(new_n1109), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n701), .B1(G50), .B2(new_n1049), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n747), .A2(new_n1055), .B1(new_n733), .B2(new_n796), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n744), .A2(G137), .ZN(new_n1127));
  INV_X1    g0927(.A(G128), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n741), .C1(new_n735), .C2(new_n1054), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1126), .B(new_n1129), .C1(G150), .C2(new_n738), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1133));
  AOI211_X1 g0933(.A(G33), .B(G41), .C1(new_n724), .C2(G124), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n788), .B2(new_n728), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT115), .Z(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1067), .A2(G58), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT114), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n742), .A2(G107), .B1(new_n746), .B2(G116), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n752), .C2(new_n723), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n283), .B(new_n396), .C1(new_n735), .C2(new_n234), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n733), .A2(new_n205), .B1(new_n743), .B2(new_n262), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1141), .A2(new_n913), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT58), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1144), .A2(KEYINPUT58), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n202), .B1(new_n381), .B2(G41), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1137), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1125), .B1(new_n1148), .B2(new_n710), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1122), .A2(new_n699), .B1(new_n1124), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1094), .A2(new_n1082), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT57), .B1(new_n1151), .B2(new_n1122), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1091), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT57), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n700), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1150), .B1(new_n1152), .B2(new_n1155), .ZN(G375));
  NAND3_X1  g0956(.A1(new_n1091), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT118), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1091), .A2(KEYINPUT118), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1159), .A2(new_n959), .A3(new_n1096), .A4(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n742), .A2(G283), .B1(new_n746), .B2(G294), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n396), .C1(new_n348), .C2(new_n728), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n733), .A2(new_n573), .B1(new_n723), .B2(new_n564), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n735), .A2(new_n205), .B1(new_n743), .B2(new_n206), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1163), .A2(new_n993), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n396), .B1(new_n744), .B2(G150), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1139), .B(new_n1167), .C1(new_n202), .C2(new_n912), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n747), .A2(new_n796), .B1(new_n741), .B2(new_n916), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n733), .A2(new_n1054), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1168), .B1(KEYINPUT119), .B2(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n735), .A2(new_n788), .B1(new_n723), .B2(new_n1128), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT120), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n1171), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1166), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n701), .B1(G68), .B2(new_n1049), .C1(new_n1178), .C2(new_n762), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n816), .B2(new_n705), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1087), .B2(new_n699), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1161), .A2(new_n1181), .ZN(G381));
  OR2_X1    g0982(.A1(G375), .A2(G378), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G393), .A2(G396), .ZN(new_n1184));
  INV_X1    g0984(.A(G384), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n1011), .A4(new_n1034), .ZN(new_n1186));
  OR4_X1    g0986(.A1(G387), .A2(new_n1183), .A3(G381), .A4(new_n1186), .ZN(G407));
  OAI211_X1 g0987(.A(G407), .B(G213), .C1(G343), .C2(new_n1183), .ZN(G409));
  INV_X1    g0988(.A(KEYINPUT126), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n704), .A2(new_n765), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n978), .B2(new_n1008), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1184), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(G390), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1011), .B(new_n1034), .C1(new_n1184), .C2(new_n1191), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT124), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT101), .B1(new_n958), .B2(new_n959), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n927), .B(new_n952), .C1(new_n957), .C2(new_n693), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n698), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n973), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1196), .B1(new_n1200), .B2(new_n926), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n926), .ZN(new_n1202));
  AOI211_X1 g1002(.A(KEYINPUT124), .B(new_n1202), .C1(new_n1199), .C2(new_n973), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1195), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(G387), .A2(KEYINPUT124), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1196), .A3(new_n926), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(G378), .B(new_n1150), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT117), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT117), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1212), .A2(new_n1153), .A3(new_n952), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1118), .B2(new_n698), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1098), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT121), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n634), .A2(G213), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1157), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n654), .B1(new_n1222), .B2(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G384), .B1(new_n1224), .B2(new_n1181), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1181), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1185), .B(new_n1226), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT121), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1209), .A2(new_n1216), .A3(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1218), .A2(new_n1219), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1225), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1227), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n1232), .ZN(new_n1237));
  AND4_X1   g1037(.A1(KEYINPUT125), .A2(new_n1217), .A3(new_n1219), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1219), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1209), .B2(new_n1216), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT125), .B1(new_n1240), .B2(new_n1237), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1233), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1234), .A2(new_n1235), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT122), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G2897), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1219), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1228), .B2(new_n1245), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1244), .B1(new_n1255), .B2(new_n1240), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1208), .B1(new_n1243), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT63), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1236), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1217), .A2(new_n1219), .A3(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1204), .A2(new_n1207), .A3(new_n1244), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1231), .B2(new_n1259), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1253), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1230), .A2(new_n1219), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1229), .B1(new_n1209), .B2(new_n1216), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT123), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1270), .B(new_n1265), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1264), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1189), .B1(new_n1258), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1264), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1256), .B1(new_n1233), .B2(new_n1242), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1274), .B(KEYINPUT126), .C1(new_n1275), .C2(new_n1208), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(G405));
  XNOR2_X1  g1077(.A(G375), .B(new_n1098), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(new_n1236), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(new_n1208), .ZN(G402));
endmodule


