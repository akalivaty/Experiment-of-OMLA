//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n541, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n470), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n466), .B1(new_n474), .B2(G2105), .ZN(G160));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n462), .A2(new_n491), .A3(G138), .A4(new_n463), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(G164));
  XNOR2_X1  g068(.A(KEYINPUT5), .B(G543), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n494), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT6), .B(G651), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n498), .A3(G88), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(G50), .A3(G543), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT69), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT69), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(G303));
  INV_X1    g078(.A(G303), .ZN(G166));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n505));
  NAND3_X1  g080(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n494), .A2(G63), .A3(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n498), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G51), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n496), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n511), .A2(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n510), .A2(new_n522), .ZN(G168));
  AOI22_X1  g098(.A1(new_n494), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n496), .B1(new_n524), .B2(KEYINPUT71), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n525), .B1(KEYINPUT71), .B2(new_n524), .ZN(new_n526));
  INV_X1    g101(.A(new_n520), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n517), .A2(new_n519), .A3(G543), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(G90), .B1(new_n528), .B2(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  NAND4_X1  g106(.A1(new_n517), .A2(new_n519), .A3(G43), .A4(G543), .ZN(new_n532));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(new_n516), .A3(G56), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n496), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT72), .Z(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G188));
  NAND3_X1  g120(.A1(new_n514), .A2(new_n516), .A3(G65), .ZN(new_n546));
  NAND2_X1  g121(.A1(G78), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(G91), .A2(new_n527), .B1(new_n548), .B2(G651), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n517), .A2(new_n519), .A3(G53), .A4(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n498), .A2(new_n552), .A3(G53), .A4(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(G299));
  INV_X1    g130(.A(G168), .ZN(G286));
  NAND2_X1  g131(.A1(new_n527), .A2(G87), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n528), .A2(G49), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n494), .B2(G74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(G288));
  AOI22_X1  g135(.A1(new_n527), .A2(G86), .B1(new_n528), .B2(G48), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n514), .A2(new_n516), .A3(G61), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n494), .A2(new_n564), .A3(G61), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n567), .A2(new_n568), .A3(G651), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n568), .B1(new_n567), .B2(G651), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n561), .B1(new_n569), .B2(new_n570), .ZN(G305));
  XNOR2_X1  g146(.A(KEYINPUT75), .B(G85), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n494), .A2(new_n498), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G47), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n494), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n573), .B1(new_n511), .B2(new_n574), .C1(new_n575), .C2(new_n496), .ZN(G290));
  INV_X1    g151(.A(G868), .ZN(new_n577));
  NOR2_X1   g152(.A1(G171), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n579));
  INV_X1    g154(.A(G92), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n520), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n494), .A2(new_n498), .A3(KEYINPUT10), .A4(G92), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n514), .A2(new_n516), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(new_n528), .B2(G54), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(G868), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT76), .B1(new_n578), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(KEYINPUT76), .B2(new_n578), .ZN(G284));
  OAI21_X1  g168(.A(new_n592), .B1(KEYINPUT76), .B2(new_n578), .ZN(G321));
  NAND2_X1  g169(.A1(G299), .A2(new_n577), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n577), .B2(G168), .ZN(G280));
  XNOR2_X1  g171(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(new_n598), .B2(G860), .ZN(G148));
  NAND2_X1  g174(.A1(new_n590), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n538), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g178(.A1(new_n477), .A2(G123), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n479), .A2(G135), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n463), .A2(G111), .ZN(new_n606));
  OAI21_X1  g181(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2096), .Z(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(G2100), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n611), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(G2443), .B(G2446), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2430), .ZN(new_n620));
  INV_X1    g195(.A(G2435), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2430), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(KEYINPUT15), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT15), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G2430), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n624), .A2(new_n626), .A3(new_n621), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n619), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n626), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2435), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n620), .A2(new_n621), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(new_n618), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT80), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n628), .A2(new_n635), .A3(new_n632), .A4(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n637), .B1(new_n634), .B2(new_n636), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n634), .A2(new_n636), .ZN(new_n644));
  INV_X1    g219(.A(new_n637), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n646), .B2(new_n638), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n617), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n641), .B1(new_n639), .B2(new_n640), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n643), .A3(new_n638), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(new_n616), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(G14), .ZN(new_n655));
  INV_X1    g230(.A(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n616), .B1(new_n651), .B2(new_n652), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n649), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n650), .B1(new_n648), .B2(new_n653), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT81), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(KEYINPUT17), .A3(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n669), .B(new_n670), .C1(new_n671), .C2(new_n668), .ZN(new_n672));
  INV_X1    g247(.A(new_n668), .ZN(new_n673));
  OAI21_X1  g248(.A(KEYINPUT18), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT82), .B(G2096), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n685), .A2(new_n686), .ZN(new_n696));
  INV_X1    g271(.A(new_n687), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(new_n691), .A3(new_n688), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n687), .B1(new_n685), .B2(new_n686), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n693), .B1(new_n688), .B2(new_n691), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n695), .A2(new_n699), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT85), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n688), .A2(new_n691), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n705), .A2(new_n694), .B1(new_n692), .B2(new_n700), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT85), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n706), .A2(new_n707), .A3(new_n702), .A4(new_n699), .ZN(new_n708));
  INV_X1    g283(.A(G1991), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n682), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n704), .A2(new_n708), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G1991), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n714), .A2(G1996), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n712), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n712), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n681), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n712), .A2(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(new_n717), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n712), .A2(new_n716), .A3(new_n718), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n723), .A2(new_n680), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(G229));
  INV_X1    g301(.A(KEYINPUT97), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n727), .A2(G2072), .B1(G29), .B2(G33), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n460), .A2(G103), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT95), .B(KEYINPUT25), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n462), .A2(G139), .A3(new_n463), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n462), .A2(G127), .ZN(new_n735));
  NAND2_X1  g310(.A1(G115), .A2(G2104), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n463), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n728), .B1(new_n738), .B2(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n727), .A2(G2072), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n739), .B(new_n740), .Z(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n490), .A2(new_n492), .ZN(new_n743));
  INV_X1    g318(.A(new_n488), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT86), .B(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G27), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n741), .B1(new_n742), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n462), .A2(G140), .A3(new_n463), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n477), .A2(G128), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n748), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  INV_X1    g337(.A(new_n750), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(G2078), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G299), .ZN(new_n765));
  INV_X1    g340(.A(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT23), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(G20), .ZN(new_n768));
  MUX2_X1   g343(.A(KEYINPUT23), .B(new_n767), .S(new_n768), .Z(new_n769));
  OAI211_X1 g344(.A(new_n751), .B(new_n764), .C1(G1956), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G1956), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n766), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n766), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT99), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT24), .B(G34), .ZN(new_n776));
  AOI22_X1  g351(.A1(G160), .A2(G29), .B1(new_n748), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  OAI22_X1  g353(.A1(new_n774), .A2(new_n775), .B1(new_n778), .B2(G2084), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n775), .B2(new_n774), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n748), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n748), .ZN(new_n782));
  MUX2_X1   g357(.A(new_n781), .B(new_n782), .S(KEYINPUT100), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2090), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n766), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n766), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G32), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT26), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n462), .A2(G129), .A3(G2105), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n462), .A2(G141), .A3(new_n463), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n460), .A2(G105), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n791), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n790), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT30), .B(G28), .Z(new_n804));
  OAI221_X1 g379(.A(new_n803), .B1(G29), .B2(new_n804), .C1(new_n608), .C2(new_n748), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT98), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n766), .A2(G19), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n538), .B2(new_n766), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1341), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n766), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n590), .B2(new_n766), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT94), .B(G1348), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n806), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  AOI211_X1 g389(.A(new_n802), .B(new_n814), .C1(G2084), .C2(new_n778), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n771), .A2(new_n780), .A3(new_n786), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n766), .A2(G22), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT91), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G166), .B2(new_n766), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT92), .B(G1971), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G16), .A2(G23), .ZN(new_n822));
  INV_X1    g397(.A(G288), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G16), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT33), .B(G1976), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  MUX2_X1   g402(.A(G6), .B(G305), .S(G16), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT32), .B(G1981), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT90), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n575), .A2(new_n496), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n573), .B1(new_n574), .B2(new_n511), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT88), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(KEYINPUT88), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(G16), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G24), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(G16), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT89), .B(G1986), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n748), .A2(G25), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n462), .A2(G131), .A3(new_n463), .ZN(new_n846));
  OR2_X1    g421(.A1(G95), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n462), .A2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(G119), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT87), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n477), .A2(G119), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT87), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n846), .A4(new_n848), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n845), .B1(new_n856), .B2(new_n748), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT35), .B(G1991), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n844), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT34), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n827), .A2(new_n861), .A3(new_n831), .A4(new_n832), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(KEYINPUT93), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(KEYINPUT93), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n834), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT36), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(new_n834), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n816), .B1(new_n867), .B2(new_n869), .ZN(G311));
  INV_X1    g445(.A(G311), .ZN(G150));
  NAND2_X1  g446(.A1(new_n535), .A2(new_n536), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G651), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n494), .A2(new_n498), .A3(G81), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n532), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT104), .B1(new_n534), .B2(new_n537), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(G55), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n527), .A2(G93), .B1(new_n528), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n494), .A2(G67), .ZN(new_n881));
  NAND2_X1  g456(.A1(G80), .A2(G543), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(G651), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT102), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G67), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n882), .B1(new_n585), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(G651), .A3(new_n883), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(new_n876), .A3(new_n877), .A4(new_n880), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n590), .A2(G559), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g473(.A(G860), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n886), .A2(G860), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT37), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(G145));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n745), .B(new_n797), .ZN(new_n905));
  INV_X1    g480(.A(new_n734), .ZN(new_n906));
  INV_X1    g481(.A(new_n737), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n757), .A3(new_n907), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n756), .B(new_n755), .C1(new_n734), .C2(new_n737), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n798), .A2(new_n745), .ZN(new_n912));
  NOR2_X1   g487(.A1(G164), .A2(new_n797), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n909), .B(new_n908), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n852), .A2(new_n855), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n462), .A2(G130), .A3(G2105), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n463), .B2(G118), .ZN(new_n920));
  INV_X1    g495(.A(G118), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(KEYINPUT105), .A3(G2105), .ZN(new_n922));
  OR2_X1    g497(.A1(G106), .A2(G2105), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n922), .A3(new_n923), .A4(G2104), .ZN(new_n924));
  INV_X1    g499(.A(G142), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n918), .B(new_n924), .C1(new_n464), .C2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n613), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n479), .A2(G142), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n613), .A3(new_n924), .A4(new_n918), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n917), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n917), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n916), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n856), .A2(new_n928), .A3(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n917), .A2(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT106), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n915), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT106), .B1(new_n935), .B2(new_n936), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n911), .A3(new_n914), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(G160), .B(new_n608), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(G162), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n904), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n941), .B2(new_n944), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(new_n938), .A3(new_n940), .A4(KEYINPUT107), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(G395));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n567), .A2(G651), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT74), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n567), .A2(new_n568), .A3(G651), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G288), .B1(new_n955), .B2(new_n561), .ZN(new_n956));
  OAI211_X1 g531(.A(G288), .B(new_n561), .C1(new_n569), .C2(new_n570), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G303), .A2(new_n837), .ZN(new_n959));
  OAI211_X1 g534(.A(G290), .B(new_n497), .C1(new_n502), .C2(new_n501), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n956), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G305), .A2(new_n823), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n963), .A2(new_n957), .B1(new_n960), .B2(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n951), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n956), .B2(new_n958), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n960), .A3(new_n959), .A4(new_n957), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(KEYINPUT110), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n894), .B(new_n600), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n548), .A2(G651), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n494), .A2(new_n498), .A3(G91), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n554), .A2(new_n972), .A3(KEYINPUT109), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(new_n583), .A3(new_n588), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n549), .B2(new_n554), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  AND3_X1   g553(.A1(G299), .A2(new_n589), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n971), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT41), .B1(new_n977), .B2(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(G299), .A2(new_n978), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(new_n590), .A3(new_n974), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT41), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n975), .A2(new_n976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n982), .B1(new_n971), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n962), .B2(new_n964), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n970), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n970), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(G868), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n886), .A2(new_n577), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(G295));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n996), .ZN(G331));
  AND4_X1   g573(.A1(new_n892), .A2(new_n876), .A3(new_n877), .A4(new_n880), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n877), .A2(new_n876), .B1(new_n892), .B2(new_n880), .ZN(new_n1000));
  OAI21_X1  g575(.A(G171), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n887), .A2(G301), .A3(new_n893), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(G168), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G168), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n980), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n887), .A2(G301), .A3(new_n893), .ZN(new_n1006));
  AOI21_X1  g581(.A(G301), .B1(new_n887), .B2(new_n893), .ZN(new_n1007));
  OAI21_X1  g582(.A(G286), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(G168), .A3(new_n1002), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n989), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1005), .A2(new_n968), .A3(new_n965), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1008), .A2(new_n989), .A3(new_n1009), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n981), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1014));
  INV_X1    g589(.A(new_n968), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT110), .B1(new_n966), .B2(new_n967), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1013), .A2(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G37), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1012), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(KEYINPUT111), .A3(new_n1018), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n983), .A2(new_n988), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n980), .A2(KEYINPUT112), .A3(new_n986), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1027), .A2(new_n1008), .A3(new_n1028), .A4(new_n1009), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1005), .A2(new_n1029), .B1(new_n965), .B2(new_n968), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1024), .A2(new_n1025), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT44), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1024), .A2(KEYINPUT43), .A3(new_n1030), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1005), .A2(new_n1010), .B1(new_n965), .B2(new_n968), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1020), .B1(new_n1034), .B2(G37), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n1022), .A3(new_n1011), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1036), .B2(KEYINPUT43), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1032), .B1(KEYINPUT44), .B2(new_n1037), .ZN(G397));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  INV_X1    g614(.A(G40), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1040), .B(new_n466), .C1(new_n474), .C2(G2105), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(G164), .B2(G1384), .ZN(new_n1043));
  INV_X1    g618(.A(G1384), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n789), .ZN(new_n1047));
  INV_X1    g622(.A(G2084), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n745), .A2(new_n1049), .A3(new_n1044), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1041), .A2(new_n1048), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1039), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT116), .B(G8), .Z(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G168), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(KEYINPUT51), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT123), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1041), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1063), .A2(new_n1048), .B1(new_n1046), .B2(new_n789), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1062), .B(new_n1059), .C1(new_n1064), .C2(new_n1055), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1064), .A2(G168), .A3(new_n1055), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G303), .A2(G8), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT55), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1041), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT115), .B(G2090), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1045), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1043), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n745), .A2(new_n1044), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1074), .A3(new_n1042), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1078), .A3(new_n1041), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT114), .B(G1971), .Z(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1073), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1070), .B1(new_n1082), .B2(new_n1055), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1070), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G160), .A2(G40), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n1075), .B2(new_n1043), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1080), .B1(new_n1086), .B2(new_n1078), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1084), .B(G8), .C1(new_n1087), .C2(new_n1073), .ZN(new_n1088));
  NAND4_X1  g663(.A1(G160), .A2(G40), .A3(new_n1044), .A4(new_n745), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n823), .A2(G1976), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1054), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  INV_X1    g667(.A(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(new_n1054), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n952), .A2(new_n561), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G1981), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(G305), .B2(G1981), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT49), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT49), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n1098), .C1(G305), .C2(G1981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1089), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1055), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1096), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1083), .A2(new_n1088), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1076), .A2(new_n742), .A3(new_n1078), .A4(new_n1041), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1046), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(G2078), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1112), .A2(new_n1113), .B1(new_n1071), .B2(new_n775), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1111), .A2(G301), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(G301), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT124), .B(new_n1108), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1068), .A2(new_n1107), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1116), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1111), .A2(G301), .A3(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1108), .B1(new_n1121), .B2(KEYINPUT124), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n549), .A2(KEYINPUT119), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1124), .A2(KEYINPUT57), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(new_n765), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT120), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1076), .A2(new_n1078), .A3(new_n1041), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1071), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1126), .A3(new_n1132), .ZN(new_n1136));
  INV_X1    g711(.A(G2067), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1104), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1071), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(new_n589), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1135), .B1(new_n1136), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(KEYINPUT60), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1148), .B2(new_n590), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1150), .A2(KEYINPUT122), .A3(new_n589), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1145), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1134), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1146), .A3(new_n590), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT122), .B1(new_n1150), .B2(new_n589), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT60), .A4(new_n1142), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1152), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1089), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1079), .A2(G1996), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n538), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(KEYINPUT59), .B(new_n538), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1133), .B(new_n1126), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1165), .B(new_n1166), .C1(new_n1167), .C2(KEYINPUT61), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1144), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1123), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n823), .A2(new_n1093), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT117), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1103), .A2(new_n1172), .B1(G1981), .B2(G305), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1105), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1106), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1088), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1066), .A2(new_n1177), .A3(new_n1067), .ZN(new_n1178));
  AND4_X1   g753(.A1(new_n1083), .A2(new_n1106), .A3(new_n1116), .A4(new_n1088), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1068), .A2(KEYINPUT62), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1176), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  OAI21_X1  g758(.A(G8), .B1(new_n1087), .B2(new_n1073), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1184), .B2(new_n1070), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1064), .A2(G286), .A3(new_n1055), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1185), .A2(new_n1088), .A3(new_n1106), .A4(new_n1186), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1083), .A2(new_n1106), .A3(new_n1088), .A4(new_n1186), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT118), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1187), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1170), .A2(new_n1182), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1085), .A2(new_n1043), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n757), .B(new_n1137), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n797), .B(new_n682), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n917), .A2(new_n858), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n917), .A2(new_n858), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(G290), .B(G1986), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1194), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1193), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(G290), .A2(G1986), .ZN(new_n1205));
  AOI21_X1  g780(.A(KEYINPUT48), .B1(new_n1194), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1194), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT48), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1205), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1206), .B(new_n1210), .C1(new_n1194), .C2(new_n1201), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1212), .A2(KEYINPUT46), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1212), .A2(KEYINPUT46), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1207), .A2(G1996), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g790(.A(new_n1195), .B(new_n798), .C1(G1996), .C2(new_n1213), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1194), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1218), .B(KEYINPUT47), .Z(new_n1219));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1197), .B1(new_n1220), .B2(new_n1199), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1200), .A2(KEYINPUT125), .ZN(new_n1222));
  OAI22_X1  g797(.A1(new_n1221), .A2(new_n1222), .B1(G2067), .B2(new_n757), .ZN(new_n1223));
  AOI211_X1 g798(.A(new_n1211), .B(new_n1219), .C1(new_n1194), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1204), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g800(.A1(G227), .A2(new_n457), .ZN(new_n1227));
  OAI211_X1 g801(.A(G14), .B(new_n654), .C1(new_n661), .C2(KEYINPUT81), .ZN(new_n1228));
  NOR2_X1   g802(.A1(new_n658), .A2(new_n659), .ZN(new_n1229));
  OAI211_X1 g803(.A(new_n948), .B(new_n1227), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g804(.A1(G229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g805(.A(new_n1025), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1232));
  OAI211_X1 g806(.A(KEYINPUT127), .B(new_n1231), .C1(new_n1232), .C2(new_n1033), .ZN(new_n1233));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1234));
  AND2_X1   g808(.A1(new_n948), .A2(new_n1227), .ZN(new_n1235));
  NAND4_X1  g809(.A1(new_n1235), .A2(new_n663), .A3(new_n725), .A4(new_n721), .ZN(new_n1236));
  OAI21_X1  g810(.A(new_n1234), .B1(new_n1037), .B2(new_n1236), .ZN(new_n1237));
  AND2_X1   g811(.A1(new_n1233), .A2(new_n1237), .ZN(G308));
  NAND2_X1  g812(.A1(new_n1233), .A2(new_n1237), .ZN(G225));
endmodule


