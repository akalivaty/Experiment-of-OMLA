//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(new_n203), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(KEYINPUT65), .A2(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(KEYINPUT65), .A2(G68), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n216), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT68), .A4(new_n216), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n260), .A2(G77), .B1(new_n261), .B2(G50), .ZN(new_n262));
  INV_X1    g0062(.A(new_n222), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n217), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT11), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n217), .A3(G1), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n255), .B2(new_n256), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G68), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT77), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT12), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n269), .A2(new_n275), .A3(new_n203), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n277));
  INV_X1    g0077(.A(new_n269), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT12), .B1(new_n263), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n273), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n274), .B1(new_n273), .B2(new_n281), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n267), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G232), .A3(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT74), .ZN(new_n297));
  AND2_X1   g0097(.A1(G1), .A2(G13), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n259), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n295), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n296), .A2(new_n297), .B1(new_n301), .B2(G238), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(G274), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT74), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT13), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT75), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n293), .A2(new_n302), .A3(new_n308), .A4(new_n304), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(G200), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(G190), .A3(new_n309), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n284), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(G169), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n310), .A2(new_n317), .A3(G169), .A4(new_n311), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n306), .A2(G179), .A3(new_n309), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n284), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n285), .A2(G232), .A3(new_n288), .ZN(new_n323));
  INV_X1    g0123(.A(G107), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n285), .A2(G1698), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n323), .B1(new_n324), .B2(new_n285), .C1(new_n325), .C2(new_n223), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n292), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n300), .A2(new_n295), .ZN(new_n328));
  INV_X1    g0128(.A(G244), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n296), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(G190), .A3(new_n331), .ZN(new_n332));
  AOI211_X1 g0132(.A(new_n296), .B(new_n330), .C1(new_n326), .C2(new_n292), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT15), .B(G87), .Z(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n260), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  INV_X1    g0140(.A(new_n261), .ZN(new_n341));
  INV_X1    g0141(.A(G77), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n340), .A2(new_n341), .B1(new_n217), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n258), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n270), .A2(G77), .A3(new_n272), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(new_n342), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT70), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n335), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n333), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n327), .A2(new_n331), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  AND4_X1   g0155(.A1(new_n314), .A2(new_n322), .A3(new_n349), .A4(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n261), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT69), .ZN(new_n359));
  MUX2_X1   g0159(.A(new_n358), .B(new_n340), .S(new_n359), .Z(new_n360));
  OAI21_X1  g0160(.A(new_n357), .B1(new_n360), .B2(new_n338), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n258), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n270), .A2(G50), .A3(new_n272), .ZN(new_n363));
  INV_X1    g0163(.A(G50), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n269), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n285), .A2(G222), .A3(new_n288), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G33), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G77), .ZN(new_n372));
  INV_X1    g0172(.A(G223), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n367), .B(new_n372), .C1(new_n325), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n292), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n296), .B1(G226), .B2(new_n301), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n353), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n350), .A3(new_n376), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n366), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n375), .A2(KEYINPUT71), .A3(G190), .A4(new_n376), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n366), .A2(KEYINPUT9), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT9), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n362), .A2(new_n388), .A3(new_n363), .A4(new_n365), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n377), .A2(G200), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n390), .B2(KEYINPUT73), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT10), .B1(new_n377), .B2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT72), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n381), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  OAI21_X1  g0203(.A(G58), .B1(new_n220), .B2(new_n221), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n213), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n285), .B2(G20), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n369), .A2(G33), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT7), .B(new_n217), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n222), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT79), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI211_X1 g0214(.A(KEYINPUT79), .B(new_n222), .C1(new_n408), .C2(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n403), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT80), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(KEYINPUT80), .B(new_n403), .C1(new_n414), .C2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(new_n411), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n420), .A2(KEYINPUT78), .A3(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT78), .B1(new_n420), .B2(G68), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT16), .B(new_n406), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n418), .A2(new_n258), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n360), .B1(new_n271), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n270), .B1(new_n360), .B2(new_n269), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(KEYINPUT81), .A3(new_n426), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n432), .B1(new_n325), .B2(new_n290), .C1(new_n373), .C2(new_n289), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n292), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT82), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n301), .A2(new_n435), .A3(G232), .ZN(new_n436));
  INV_X1    g0236(.A(G232), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT82), .B1(new_n328), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n296), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n434), .A2(new_n439), .A3(G179), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n353), .B1(new_n434), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n429), .A2(new_n430), .A3(new_n431), .A4(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n334), .B1(new_n434), .B2(new_n439), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n434), .A2(new_n439), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n445), .B1(G190), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n424), .A2(new_n426), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n424), .A2(new_n447), .A3(KEYINPUT17), .A4(new_n426), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n429), .A2(new_n431), .A3(new_n443), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(KEYINPUT18), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n356), .A2(new_n402), .A3(new_n444), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n324), .A2(KEYINPUT6), .A3(G97), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n324), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n206), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n456), .B1(new_n459), .B2(KEYINPUT6), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n420), .A2(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n463), .A2(new_n258), .B1(new_n457), .B2(new_n269), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n271), .A2(G33), .ZN(new_n465));
  AND3_X1   g0265(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n298), .B1(new_n466), .B2(new_n251), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT68), .B1(new_n467), .B2(new_n250), .ZN(new_n468));
  INV_X1    g0268(.A(new_n256), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n278), .B(new_n465), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n270), .A2(KEYINPUT83), .A3(new_n465), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(G97), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n271), .B(G45), .C1(new_n299), .C2(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT85), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n476), .B2(KEYINPUT85), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(new_n300), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n476), .A2(KEYINPUT85), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n292), .A2(new_n294), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n477), .A4(new_n479), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n368), .A2(new_n370), .A3(G250), .A4(G1698), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT84), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n368), .A2(new_n370), .A3(G244), .A4(new_n288), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n292), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n353), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n486), .A2(new_n495), .A3(new_n350), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n475), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(G200), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n486), .A2(new_n495), .A3(G190), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(new_n464), .A3(new_n501), .A4(new_n474), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n285), .A2(G238), .A3(new_n288), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  OAI221_X1 g0305(.A(new_n504), .B1(new_n259), .B2(new_n505), .C1(new_n325), .C2(new_n329), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n292), .ZN(new_n507));
  INV_X1    g0307(.A(G45), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G1), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n294), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n300), .B(new_n510), .C1(G250), .C2(new_n509), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G179), .ZN(new_n513));
  AOI21_X1  g0313(.A(G169), .B1(new_n507), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n472), .A2(new_n336), .A3(new_n473), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n338), .B2(new_n457), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n285), .A2(new_n217), .A3(G68), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n217), .B1(new_n287), .B2(new_n518), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G87), .B2(new_n207), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n258), .A2(new_n523), .B1(new_n269), .B2(new_n337), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n517), .B1(new_n516), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n515), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n472), .A2(G87), .A3(new_n473), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n528), .A2(new_n524), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n512), .A2(G200), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n530), .C1(new_n383), .C2(new_n512), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n269), .A2(new_n324), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n532), .B(KEYINPUT25), .ZN(new_n533));
  OR3_X1    g0333(.A1(new_n217), .A2(KEYINPUT23), .A3(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n217), .A2(G33), .A3(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT23), .B1(new_n217), .B2(G107), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n285), .A2(new_n217), .A3(G87), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT91), .B(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n285), .A2(new_n540), .A3(new_n217), .A4(G87), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n257), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n533), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n285), .A2(G257), .A3(G1698), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n285), .A2(G250), .A3(new_n288), .ZN(new_n551));
  INV_X1    g0351(.A(G294), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n259), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n292), .ZN(new_n554));
  OAI211_X1 g0354(.A(G264), .B(new_n300), .C1(new_n478), .C2(new_n480), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(G190), .A3(new_n484), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n472), .A2(G107), .A3(new_n473), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n484), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n549), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n503), .A2(new_n527), .A3(new_n531), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(G20), .B1(G33), .B2(G283), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n259), .A2(G97), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(G20), .B2(new_n505), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT20), .B1(new_n253), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n253), .A2(new_n565), .A3(KEYINPUT20), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(KEYINPUT88), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n253), .A2(new_n565), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n568), .A2(new_n572), .B1(G116), .B2(new_n278), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT87), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n470), .B2(new_n505), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n270), .A2(KEYINPUT87), .A3(G116), .A4(new_n465), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n285), .A2(G257), .A3(new_n288), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n285), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n292), .ZN(new_n583));
  OAI211_X1 g0383(.A(G270), .B(new_n300), .C1(new_n478), .C2(new_n480), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n484), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n577), .A2(new_n578), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n575), .A2(new_n576), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n567), .A2(KEYINPUT88), .ZN(new_n589));
  INV_X1    g0389(.A(new_n566), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(new_n571), .B1(new_n505), .B2(new_n269), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n586), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT21), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n585), .A2(new_n350), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT89), .B1(new_n577), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT89), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n583), .A2(G190), .A3(new_n484), .A4(new_n584), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(G200), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n577), .A2(KEYINPUT90), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT90), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n603), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n593), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n549), .A2(new_n558), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n559), .A2(new_n353), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(G179), .C2(new_n559), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n596), .A2(new_n602), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n455), .A2(new_n562), .A3(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n455), .ZN(new_n615));
  INV_X1    g0415(.A(new_n499), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n527), .A2(new_n531), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n618));
  XNOR2_X1  g0418(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n527), .A2(new_n531), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n527), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT94), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT94), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n618), .A2(new_n623), .A3(new_n527), .A4(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n527), .A2(new_n531), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n499), .A2(new_n561), .A3(new_n502), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n596), .A2(new_n602), .A3(new_n612), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n622), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n615), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT95), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n351), .A2(new_n348), .A3(new_n354), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n314), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n452), .B1(new_n322), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n427), .A2(new_n443), .ZN(new_n636));
  XNOR2_X1  g0436(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n442), .B1(new_n424), .B2(new_n426), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n395), .B2(new_n401), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n381), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n632), .A2(new_n645), .ZN(G369));
  NAND2_X1  g0446(.A1(new_n596), .A2(new_n602), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n271), .A2(new_n217), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n593), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n653), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n609), .B1(new_n577), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n647), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n610), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n561), .B1(new_n659), .B2(new_n655), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n612), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n611), .B1(G179), .B2(new_n559), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n655), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n653), .B1(new_n596), .B2(new_n602), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n661), .B1(new_n663), .B2(new_n655), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n210), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n214), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(new_n619), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n617), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n527), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n627), .B2(new_n628), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n653), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n621), .A2(KEYINPUT94), .B1(new_n627), .B2(new_n628), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n653), .B1(new_n686), .B2(new_n624), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n687), .B2(KEYINPUT29), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n596), .A2(new_n602), .A3(new_n612), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n627), .A3(new_n609), .A4(new_n655), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n495), .A2(new_n484), .A3(new_n481), .ZN(new_n692));
  INV_X1    g0492(.A(new_n512), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n597), .A3(new_n693), .A4(new_n556), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n693), .A2(G179), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(new_n496), .A3(new_n559), .A4(new_n585), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n556), .A2(new_n507), .A3(new_n511), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n597), .A3(KEYINPUT30), .A4(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n691), .B1(new_n701), .B2(new_n653), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n691), .A3(new_n653), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n690), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n688), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n677), .B1(new_n709), .B2(G1), .ZN(G364));
  NOR2_X1   g0510(.A1(new_n657), .A2(G330), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT97), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n268), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n271), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n712), .B(new_n658), .C1(new_n672), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n672), .A2(new_n715), .ZN(new_n717));
  INV_X1    g0517(.A(G355), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n285), .A2(new_n210), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n718), .A2(new_n719), .B1(G116), .B2(new_n210), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n247), .A2(G45), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n671), .A2(new_n285), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n508), .B2(new_n215), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n720), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT98), .ZN(new_n726));
  OAI21_X1  g0526(.A(G20), .B1(new_n726), .B2(G169), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n353), .A2(KEYINPUT98), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n298), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT99), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n717), .B1(new_n725), .B2(new_n738), .ZN(new_n739));
  OR3_X1    g0539(.A1(new_n217), .A2(KEYINPUT100), .A3(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n334), .A2(G179), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT100), .B1(new_n217), .B2(G190), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(G283), .A2(new_n744), .B1(new_n747), .B2(G329), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n217), .A2(new_n383), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n350), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n217), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n752), .A2(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n750), .A2(new_n741), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n285), .B(new_n757), .C1(G303), .C2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n383), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n217), .B1(new_n745), .B2(G190), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n552), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n761), .A2(G190), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n749), .A2(new_n760), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n747), .A2(G159), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n759), .A2(G87), .ZN(new_n773));
  AOI21_X1  g0573(.A(KEYINPUT101), .B1(new_n773), .B2(new_n285), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G107), .B2(new_n744), .ZN(new_n775));
  INV_X1    g0575(.A(new_n767), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n776), .A2(new_n203), .B1(new_n763), .B2(new_n364), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n752), .A2(new_n202), .B1(new_n755), .B2(new_n342), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n765), .A2(new_n457), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n773), .A2(KEYINPUT101), .A3(new_n285), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n775), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n770), .B1(new_n772), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n739), .B1(new_n783), .B2(new_n733), .ZN(new_n784));
  INV_X1    g0584(.A(new_n736), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n657), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n716), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n348), .A2(new_n653), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n335), .B2(new_n348), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n355), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT104), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n633), .A2(new_n655), .ZN(new_n793));
  AND3_X1   g0593(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n655), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n686), .B2(new_n624), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n687), .B2(new_n796), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n707), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT105), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n717), .B1(new_n800), .B2(new_n707), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n733), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n735), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n717), .B1(new_n806), .B2(G77), .ZN(new_n807));
  INV_X1    g0607(.A(new_n752), .ZN(new_n808));
  INV_X1    g0608(.A(new_n755), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G143), .A2(new_n808), .B1(new_n809), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G150), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n776), .B2(new_n811), .C1(new_n812), .C2(new_n763), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n743), .A2(new_n203), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n285), .B1(new_n765), .B2(new_n202), .C1(new_n364), .C2(new_n758), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G132), .C2(new_n747), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT103), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT103), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n814), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n324), .A2(new_n758), .B1(new_n752), .B2(new_n552), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n285), .B(new_n821), .C1(G116), .C2(new_n809), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n763), .A2(new_n581), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n779), .B(new_n823), .C1(G283), .C2(new_n767), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n747), .A2(G311), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n744), .A2(G87), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n807), .B1(new_n828), .B2(new_n733), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n796), .B2(new_n735), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n804), .A2(new_n830), .ZN(G384));
  NAND2_X1  g0631(.A1(new_n642), .A2(new_n651), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT38), .ZN(new_n833));
  INV_X1    g0633(.A(new_n651), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n429), .A2(new_n431), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n448), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n453), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n424), .A2(new_n426), .A3(new_n447), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n406), .B1(new_n422), .B2(new_n421), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n403), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n258), .A3(new_n423), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n843), .A2(new_n426), .B1(new_n442), .B2(new_n651), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n453), .A2(KEYINPUT18), .ZN(new_n846));
  INV_X1    g0646(.A(new_n452), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n444), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n651), .B1(new_n843), .B2(new_n426), .ZN(new_n849));
  AOI221_X4 g0649(.A(new_n833), .B1(new_n839), .B2(new_n845), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n839), .A2(new_n845), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n321), .A2(new_n653), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n322), .A2(new_n314), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n314), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n321), .B(new_n653), .C1(new_n320), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n793), .B(KEYINPUT106), .Z(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n798), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n832), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT107), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n452), .A2(KEYINPUT109), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n640), .B(new_n638), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT109), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n450), .A2(new_n868), .A3(new_n451), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n431), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT81), .B1(new_n424), .B2(new_n426), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n871), .A2(new_n872), .A3(new_n651), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n448), .A2(KEYINPUT108), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT108), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n424), .A2(new_n447), .A3(new_n876), .A4(new_n426), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n636), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n839), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n865), .B1(new_n850), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n322), .A2(new_n653), .ZN(new_n883));
  INV_X1    g0683(.A(new_n849), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n454), .B2(new_n444), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n839), .A2(new_n845), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n833), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n882), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT107), .B(new_n832), .C1(new_n854), .C2(new_n861), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n864), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n615), .B(new_n685), .C1(new_n687), .C2(KEYINPUT29), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n645), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(G330), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n794), .A2(new_n795), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n856), .B2(new_n858), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n706), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n887), .B2(new_n888), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n706), .A2(new_n898), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n850), .B2(new_n881), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n904), .B2(KEYINPUT40), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n615), .A2(new_n706), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n905), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n895), .A2(new_n908), .B1(new_n271), .B2(new_n713), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT110), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n895), .A2(new_n908), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n915), .A2(G116), .A3(new_n218), .A4(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT36), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n215), .A2(G77), .A3(new_n404), .ZN(new_n919));
  INV_X1    g0719(.A(new_n201), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n203), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n268), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n918), .A3(new_n922), .ZN(G367));
  INV_X1    g0723(.A(new_n669), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n475), .A2(new_n653), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n503), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n616), .A2(new_n653), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT112), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT112), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n669), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n669), .A2(new_n928), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT44), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n666), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n935), .A2(new_n667), .A3(new_n938), .A4(new_n936), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n665), .B(new_n668), .Z(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n658), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n709), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n672), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n714), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT113), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT111), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n666), .B2(new_n928), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n529), .A2(new_n655), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n527), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n527), .A2(new_n954), .A3(new_n531), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n666), .A2(new_n951), .A3(new_n928), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n953), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n953), .B2(new_n960), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n928), .A2(new_n668), .A3(new_n664), .A4(new_n661), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n503), .A2(new_n663), .A3(new_n925), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n653), .B1(new_n965), .B2(new_n499), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n963), .B2(KEYINPUT42), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n964), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n961), .A2(new_n962), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n961), .B2(new_n962), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n949), .A2(new_n950), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n715), .B1(new_n945), .B2(new_n947), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT113), .B1(new_n975), .B2(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n955), .A2(new_n736), .A3(new_n956), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n239), .A2(new_n723), .B1(new_n210), .B2(new_n337), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n717), .B1(new_n738), .B2(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n752), .A2(new_n811), .B1(new_n755), .B2(new_n201), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n371), .B(new_n981), .C1(G58), .C2(new_n759), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n744), .A2(G77), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n812), .C2(new_n746), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n765), .A2(new_n203), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n762), .A2(G143), .ZN(new_n987));
  INV_X1    g0787(.A(G159), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n776), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n808), .A2(G303), .B1(G311), .B2(new_n762), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT114), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n758), .A2(new_n505), .ZN(new_n992));
  INV_X1    g0792(.A(new_n765), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n992), .A2(KEYINPUT46), .B1(G107), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(KEYINPUT114), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n992), .A2(KEYINPUT46), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n991), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n744), .A2(G97), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT115), .B(G317), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n747), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n767), .A2(G294), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n285), .B1(new_n809), .B2(G283), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n984), .A2(new_n989), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT47), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n805), .B1(new_n1005), .B2(KEYINPUT47), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n980), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n978), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n977), .A2(new_n1009), .ZN(G387));
  NOR2_X1   g0810(.A1(new_n236), .A2(new_n508), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n340), .A2(G50), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT50), .Z(new_n1013));
  OAI211_X1 g0813(.A(new_n674), .B(new_n508), .C1(new_n203), .C2(new_n342), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n722), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1011), .B1(KEYINPUT116), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT116), .B2(new_n1015), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(G107), .B2(new_n210), .C1(new_n674), .C2(new_n719), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n737), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n998), .B1(new_n811), .B2(new_n746), .C1(new_n360), .C2(new_n776), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G77), .A2(new_n759), .B1(new_n809), .B2(G68), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n285), .C1(new_n364), .C2(new_n752), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n993), .A2(new_n336), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n763), .B2(new_n988), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n808), .A2(new_n999), .B1(new_n809), .B2(G303), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n776), .B2(new_n756), .C1(new_n753), .C2(new_n763), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  INV_X1    g0830(.A(G283), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n758), .A2(new_n552), .B1(new_n765), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT117), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n371), .B1(new_n743), .B2(new_n505), .C1(new_n764), .C2(new_n746), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1025), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1019), .B(new_n717), .C1(new_n805), .C2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n665), .B2(new_n736), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n944), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n715), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n709), .A2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n672), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n709), .A2(new_n1042), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  AND2_X1   g0847(.A1(new_n940), .A2(new_n941), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1044), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n673), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n244), .A2(new_n723), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n737), .B1(new_n457), .B2(new_n210), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n717), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT118), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n763), .A2(new_n811), .B1(new_n752), .B2(new_n988), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT51), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n285), .B1(new_n755), .B2(new_n340), .C1(new_n222), .C2(new_n758), .ZN(new_n1059));
  INV_X1    g0859(.A(G143), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n826), .B1(new_n1060), .B2(new_n746), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n776), .A2(new_n201), .B1(new_n342), .B2(new_n765), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n808), .A2(G311), .B1(G317), .B2(new_n762), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n371), .B1(new_n755), .B2(new_n552), .C1(new_n1031), .C2(new_n758), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n776), .A2(new_n581), .B1(new_n765), .B2(new_n505), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n324), .A2(new_n743), .B1(new_n746), .B2(new_n753), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n733), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1056), .B(new_n1072), .C1(new_n929), .C2(new_n736), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1048), .B2(new_n715), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1051), .A2(new_n1074), .ZN(G390));
  AND3_X1   g0875(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n868), .B1(new_n450), .B2(new_n451), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n642), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n835), .B1(new_n1078), .B2(new_n869), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n871), .A2(new_n872), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n837), .B1(new_n1080), .B2(new_n443), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n448), .A2(KEYINPUT108), .B1(new_n427), .B2(new_n443), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n835), .A2(new_n877), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n835), .A2(new_n1081), .B1(new_n1083), .B2(KEYINPUT37), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n833), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT39), .B1(new_n1085), .B2(new_n888), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n734), .B1(new_n1076), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n765), .A2(new_n342), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n763), .A2(new_n1031), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G107), .C2(new_n767), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n746), .A2(new_n552), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G116), .A2(new_n808), .B1(new_n809), .B2(G97), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n371), .A3(new_n773), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1091), .A2(new_n815), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1097));
  INV_X1    g0897(.A(G132), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n285), .B1(new_n752), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n759), .A2(G150), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1100), .A2(KEYINPUT53), .B1(new_n812), .B2(new_n776), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1099), .B(new_n1101), .C1(new_n809), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(KEYINPUT53), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n993), .A2(G159), .B1(G128), .B2(new_n762), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G125), .A2(new_n747), .B1(new_n744), .B2(new_n920), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1096), .A2(new_n1097), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n733), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n805), .A2(new_n360), .A3(new_n735), .ZN(new_n1111));
  AND4_X1   g0911(.A1(new_n717), .A2(new_n1087), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n896), .B1(new_n690), .B2(new_n705), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n796), .A3(new_n859), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n883), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n882), .A2(new_n889), .B1(new_n861), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1085), .A2(new_n888), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n653), .B(new_n897), .C1(new_n681), .C2(new_n683), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n859), .B1(new_n1119), .B2(new_n860), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1118), .A2(new_n1120), .A3(new_n1116), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1115), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n797), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n860), .B1(new_n630), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n859), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1076), .B2(new_n1086), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n1114), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1112), .B1(new_n1131), .B2(new_n715), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n613), .A2(new_n562), .A3(new_n653), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n701), .A2(new_n691), .A3(new_n653), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n702), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n796), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1125), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1124), .B1(new_n1114), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n860), .B1(new_n684), .B2(new_n796), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1139), .A2(new_n1114), .A3(new_n1137), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT119), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n707), .B2(new_n455), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n356), .A2(new_n402), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n848), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n1113), .A3(KEYINPUT119), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n893), .A3(new_n645), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1122), .A2(new_n1129), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(KEYINPUT120), .A3(new_n672), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1131), .B2(new_n1149), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT120), .B1(new_n1150), .B2(new_n672), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1132), .B1(new_n1152), .B2(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n1148), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n366), .A2(new_n834), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n402), .B(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1158), .B(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n905), .A2(new_n1161), .A3(new_n896), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1158), .B(new_n1159), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n899), .B(new_n903), .C1(new_n850), .C2(new_n853), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n902), .B1(new_n1085), .B2(new_n888), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n899), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1163), .B1(new_n1166), .B2(G330), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n892), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n891), .A2(new_n890), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1161), .B1(new_n905), .B2(new_n896), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n899), .B1(new_n1118), .B2(new_n903), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1163), .B(G330), .C1(new_n1171), .C2(new_n901), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n864), .A2(new_n1169), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1156), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n673), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n892), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1169), .A2(new_n1170), .A3(new_n864), .A4(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1156), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT123), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT123), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1182), .A3(KEYINPUT57), .A4(new_n1156), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1176), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n776), .A2(new_n1098), .B1(new_n765), .B2(new_n811), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G128), .A2(new_n808), .B1(new_n759), .B2(new_n1103), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n812), .B2(new_n755), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G125), .C2(new_n762), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n259), .B(new_n299), .C1(new_n743), .C2(new_n988), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G124), .B2(new_n747), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n986), .B1(new_n776), .B2(new_n457), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n337), .A2(new_n755), .B1(new_n324), .B2(new_n752), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n299), .B(new_n371), .C1(new_n758), .C2(new_n342), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n744), .A2(G58), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n1031), .C2(new_n746), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1195), .B(new_n1200), .C1(G116), .C2(new_n762), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT58), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G50), .B1(new_n259), .B2(new_n299), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n285), .B2(G41), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1194), .A2(new_n1202), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n733), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n717), .C1(new_n920), .C2(new_n806), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1161), .B2(new_n734), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1179), .B2(new_n715), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1184), .A2(new_n1211), .ZN(G375));
  INV_X1    g1012(.A(new_n1141), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n714), .B(KEYINPUT124), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n717), .B1(new_n806), .B2(G68), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n758), .A2(new_n988), .B1(new_n755), .B2(new_n811), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n371), .B(new_n1217), .C1(G137), .C2(new_n808), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n763), .A2(new_n1098), .B1(new_n765), .B2(new_n364), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n767), .B2(new_n1103), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n747), .A2(G128), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1199), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n983), .A2(new_n371), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT125), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1023), .B1(new_n776), .B2(new_n505), .C1(new_n552), .C2(new_n763), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n758), .A2(new_n457), .B1(new_n755), .B2(new_n324), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G283), .B2(new_n808), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n581), .C2(new_n746), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1216), .B1(new_n1230), .B2(new_n733), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n859), .B2(new_n735), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1215), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n947), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1235), .B2(new_n1237), .ZN(G381));
  INV_X1    g1038(.A(G375), .ZN(new_n1239));
  INV_X1    g1039(.A(G390), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1242), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n974), .A2(new_n976), .B1(new_n978), .B2(new_n1008), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1239), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n652), .A2(G213), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(new_n1249), .C2(G375), .ZN(G409));
  XNOR2_X1  g1050(.A(G393), .B(new_n787), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1251), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1244), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1240), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1244), .B2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1257), .B(G390), .C1(new_n1244), .C2(new_n1253), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1184), .A2(G378), .A3(new_n1211), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1210), .B1(new_n1179), .B2(new_n1214), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n946), .B2(new_n1174), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1245), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1248), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1236), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n672), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1234), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1241), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G384), .A2(new_n1234), .A3(new_n1269), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1248), .A2(G2897), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1273), .B(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1260), .B1(new_n1265), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1273), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1265), .B2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1248), .B(new_n1273), .C1(new_n1261), .C2(new_n1264), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1278), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1259), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1260), .C1(new_n1265), .C2(new_n1276), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1259), .B1(new_n1282), .B2(KEYINPUT63), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT127), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1277), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1265), .A2(new_n1279), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1294), .A3(new_n1259), .A4(new_n1285), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1290), .B(new_n1295), .C1(new_n1297), .C2(new_n1259), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1289), .A2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1245), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1261), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1273), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1259), .ZN(G402));
endmodule


