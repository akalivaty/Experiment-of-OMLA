//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT74), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G141gat), .B(G148gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n204), .B(new_n210), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n220), .A2(KEYINPUT75), .A3(new_n204), .A4(new_n210), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n213), .B(KEYINPUT76), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n209), .A2(KEYINPUT77), .A3(KEYINPUT2), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n202), .A2(new_n203), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT77), .B1(new_n209), .B2(KEYINPUT2), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n222), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT29), .ZN(new_n231));
  INV_X1    g030(.A(G211gat), .ZN(new_n232));
  INV_X1    g031(.A(G218gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(G211gat), .B2(G218gat), .ZN(new_n237));
  XOR2_X1   g036(.A(G197gat), .B(G204gat), .Z(new_n238));
  OR2_X1    g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G211gat), .A2(G218gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(new_n234), .C1(new_n238), .C2(new_n235), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n231), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n216), .A2(new_n221), .B1(new_n224), .B2(new_n228), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n246), .B2(new_n223), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n241), .B(KEYINPUT79), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n239), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n251), .B2(new_n245), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n252), .B2(new_n244), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n248), .A2(new_n249), .B1(new_n253), .B2(new_n243), .ZN(new_n254));
  XOR2_X1   g053(.A(G78gat), .B(G106gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G22gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT31), .B(G50gat), .Z(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  XOR2_X1   g057(.A(new_n254), .B(new_n258), .Z(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(KEYINPUT1), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n260), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n222), .A2(new_n229), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n267), .ZN(new_n271));
  INV_X1    g070(.A(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n244), .B2(new_n223), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n270), .B(new_n271), .C1(new_n273), .C2(new_n230), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT39), .ZN(new_n275));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G57gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  AND2_X1   g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(new_n277), .ZN(new_n284));
  INV_X1    g083(.A(new_n268), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n244), .A2(new_n267), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n284), .B(KEYINPUT39), .C1(new_n287), .C2(new_n277), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT40), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n277), .B1(new_n285), .B2(new_n286), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n285), .A2(new_n276), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT5), .B(new_n291), .C1(new_n274), .C2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n273), .A2(new_n230), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n294), .A2(new_n271), .A3(new_n270), .A4(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n290), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(new_n290), .A3(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n282), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n289), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n288), .A3(KEYINPUT40), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT81), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT81), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n283), .A2(new_n288), .A3(new_n305), .A4(KEYINPUT40), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G226gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  OR2_X1    g112(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n315));
  AOI21_X1  g114(.A(G190gat), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(KEYINPUT25), .B(new_n313), .C1(new_n316), .C2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n319), .A2(new_n333), .A3(new_n320), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n312), .B2(KEYINPUT23), .ZN(new_n336));
  AND4_X1   g135(.A1(new_n335), .A2(new_n324), .A3(new_n325), .A4(KEYINPUT23), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n328), .B(new_n334), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n330), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT26), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n312), .B2(new_n345), .ZN(new_n346));
  NOR3_X1   g145(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n317), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n350), .B(new_n317), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT27), .B(G183gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(KEYINPUT28), .A3(new_n332), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n352), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n332), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n314), .A2(KEYINPUT27), .A3(new_n315), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(KEYINPUT27), .B2(G183gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n361), .B2(new_n332), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n349), .B(new_n351), .C1(new_n357), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n311), .B1(new_n343), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n343), .B2(new_n363), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n366), .A2(new_n367), .A3(new_n310), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n322), .A2(new_n329), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n338), .A2(new_n340), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT65), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n349), .A2(new_n351), .ZN(new_n374));
  INV_X1    g173(.A(new_n357), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n361), .A2(new_n332), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n358), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n245), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT71), .B1(new_n379), .B2(new_n311), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n365), .B1(new_n368), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n242), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n311), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(new_n242), .A3(new_n365), .ZN(new_n386));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  NAND4_X1  g190(.A1(new_n383), .A2(new_n384), .A3(new_n386), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n367), .B1(new_n366), .B2(new_n310), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT71), .A3(new_n311), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n242), .B1(new_n396), .B2(new_n365), .ZN(new_n397));
  INV_X1    g196(.A(new_n386), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n364), .B1(new_n394), .B2(new_n395), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n386), .B(new_n391), .C1(new_n400), .C2(new_n242), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n302), .A2(new_n307), .A3(new_n392), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n282), .B1(new_n293), .B2(new_n296), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n404), .A2(KEYINPUT82), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT82), .B1(new_n404), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n299), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n301), .B1(new_n409), .B2(new_n297), .ZN(new_n410));
  INV_X1    g209(.A(new_n405), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n293), .A2(new_n296), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n301), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n386), .B1(new_n400), .B2(new_n242), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n393), .B1(new_n416), .B2(KEYINPUT37), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT38), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n385), .A2(new_n382), .A3(new_n365), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n400), .B2(new_n382), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n408), .B(new_n415), .C1(new_n417), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n383), .B2(new_n386), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT38), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n401), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n259), .B(new_n403), .C1(new_n423), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n392), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n404), .A2(new_n405), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n413), .B2(new_n404), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n259), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n373), .A2(new_n378), .A3(new_n272), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n267), .B1(new_n343), .B2(new_n363), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n272), .B1(new_n373), .B2(new_n378), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n343), .A2(new_n267), .A3(new_n363), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n432), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(KEYINPUT33), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n432), .A3(new_n445), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT34), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT70), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n444), .A2(KEYINPUT34), .A3(new_n432), .A4(new_n445), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n443), .B(new_n450), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT70), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n447), .A2(new_n449), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n445), .ZN(new_n462));
  AOI221_X4 g261(.A(new_n448), .B1(KEYINPUT33), .B2(new_n442), .C1(new_n462), .C2(new_n433), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n431), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n427), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n408), .A2(new_n415), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n254), .B(new_n258), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n428), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n474), .A2(new_n430), .A3(new_n428), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n475), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G43gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(KEYINPUT87), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n481), .B1(new_n485), .B2(G43gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G43gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G50gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT15), .ZN(new_n495));
  NAND2_X1  g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT86), .Z(new_n497));
  NOR2_X1   g296(.A1(G29gat), .A2(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n500), .A2(G29gat), .A3(G36gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n488), .A2(new_n495), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT15), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n499), .B2(new_n501), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n498), .A2(KEYINPUT14), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT85), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n497), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n503), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n503), .B2(new_n511), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT89), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT16), .ZN(new_n519));
  OR2_X1    g318(.A1(G15gat), .A2(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g320(.A1(G15gat), .A2(G22gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G8gat), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n517), .A2(new_n523), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(G1gat), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n517), .A2(new_n519), .A3(new_n523), .ZN(new_n528));
  AOI21_X1  g327(.A(G1gat), .B1(new_n517), .B2(new_n523), .ZN(new_n529));
  OAI21_X1  g328(.A(G8gat), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n515), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT13), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n527), .A2(new_n530), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n513), .B2(new_n514), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n503), .A2(new_n511), .A3(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT91), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n515), .A2(new_n531), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n540), .A2(new_n542), .A3(new_n547), .A4(new_n543), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n545), .A2(new_n533), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n536), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(KEYINPUT92), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n554), .A3(new_n550), .ZN(new_n555));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT12), .Z(new_n561));
  AND2_X1   g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n545), .A2(new_n548), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n546), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n552), .A3(new_n536), .ZN(new_n565));
  INV_X1    g364(.A(new_n561), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n553), .A2(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(G64gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G57gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n569), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(KEYINPUT94), .A3(new_n573), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  INV_X1    g377(.A(new_n573), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n575), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n573), .B(KEYINPUT93), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n583), .A2(new_n574), .A3(new_n575), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n591), .A2(new_n592), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n597), .B2(new_n588), .ZN(new_n598));
  OAI22_X1  g397(.A1(new_n582), .A2(new_n584), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g399(.A(new_n574), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n573), .B(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n603), .A3(new_n576), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n593), .A2(new_n595), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n594), .A3(new_n588), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .A4(new_n581), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT97), .B1(new_n607), .B2(new_n600), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n582), .A2(new_n584), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n596), .A2(new_n598), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .A4(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT98), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  INV_X1    g418(.A(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(G176gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n599), .A2(new_n607), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n616), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n618), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n618), .A2(KEYINPUT101), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n629), .A3(new_n617), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n628), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n623), .B(KEYINPUT100), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n627), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n567), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n638), .A2(new_n531), .A3(G183gat), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640));
  OAI21_X1  g439(.A(G183gat), .B1(new_n638), .B2(new_n531), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n640), .B1(new_n639), .B2(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n636), .A3(new_n642), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT20), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G211gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n645), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n645), .B2(new_n647), .ZN(new_n653));
  XOR2_X1   g452(.A(G127gat), .B(G155gat), .Z(new_n654));
  NAND2_X1  g453(.A1(G231gat), .A2(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n652), .B2(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n515), .A2(new_n611), .ZN(new_n662));
  NAND3_X1  g461(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n542), .A2(new_n543), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n611), .ZN(new_n665));
  XNOR2_X1  g464(.A(G190gat), .B(G218gat), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G134gat), .B(G162gat), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n667), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n479), .A2(new_n635), .A3(new_n661), .A4(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n430), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n518), .ZN(G1324gat));
  OAI21_X1  g480(.A(G8gat), .B1(new_n679), .B2(new_n428), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  INV_X1    g482(.A(new_n428), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n525), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n684), .B(new_n686), .C1(new_n677), .C2(new_n678), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n691));
  OAI221_X1 g490(.A(new_n682), .B1(new_n683), .B2(new_n687), .C1(new_n690), .C2(new_n691), .ZN(G1325gat));
  INV_X1    g491(.A(new_n679), .ZN(new_n693));
  INV_X1    g492(.A(new_n465), .ZN(new_n694));
  AOI21_X1  g493(.A(G15gat), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n469), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(G15gat), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n679), .A2(new_n259), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n471), .A2(KEYINPUT106), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n427), .A2(new_n470), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n478), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n705), .B2(new_n674), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n675), .B1(new_n471), .B2(new_n478), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n635), .A2(new_n660), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n712), .B2(new_n430), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  INV_X1    g513(.A(new_n430), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n710), .A2(new_n714), .A3(new_n715), .A4(new_n711), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(G29gat), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n707), .A2(new_n711), .ZN(new_n718));
  INV_X1    g517(.A(G29gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n719), .A3(new_n715), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(G1328gat));
  INV_X1    g521(.A(G36gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n723), .A3(new_n684), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT46), .Z(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n712), .B2(new_n428), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n469), .A3(new_n711), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n718), .A2(new_n489), .A3(new_n694), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n705), .A2(new_n674), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n473), .A2(new_n738), .A3(new_n711), .A4(new_n708), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(new_n485), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n718), .A2(new_n485), .A3(new_n473), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n739), .B2(new_n485), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  OAI221_X1 g543(.A(new_n741), .B1(new_n735), .B2(KEYINPUT48), .C1(new_n739), .C2(new_n485), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1331gat));
  NAND2_X1  g545(.A1(new_n565), .A2(new_n566), .ZN(new_n747));
  INV_X1    g546(.A(new_n551), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n749), .A3(new_n561), .A4(new_n555), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n660), .A2(new_n674), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n705), .A2(new_n634), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n705), .A2(KEYINPUT109), .A3(new_n634), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n430), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n568), .ZN(G1332gat));
  NAND2_X1  g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n755), .A2(new_n684), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(KEYINPUT110), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(KEYINPUT110), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n755), .A2(new_n756), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(new_n768), .A3(new_n684), .A4(new_n760), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n761), .A2(KEYINPUT110), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n766), .A2(new_n771), .ZN(G1333gat));
  NAND3_X1  g571(.A1(new_n767), .A2(G71gat), .A3(new_n469), .ZN(new_n773));
  INV_X1    g572(.A(G71gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n757), .B2(new_n465), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT50), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n757), .A2(new_n259), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT111), .B(G78gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n661), .A2(new_n751), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n634), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n706), .A2(new_n709), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n430), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  INV_X1    g588(.A(new_n784), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n736), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n674), .A4(new_n784), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n715), .A2(new_n634), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n586), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT112), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n788), .B1(new_n793), .B2(new_n797), .ZN(G1336gat));
  AOI21_X1  g597(.A(new_n587), .B1(new_n786), .B2(new_n684), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n684), .A2(new_n587), .A3(new_n634), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT113), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n800), .B(new_n801), .C1(new_n793), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n793), .A2(new_n804), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n806), .B2(new_n799), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n787), .B2(new_n696), .ZN(new_n809));
  INV_X1    g608(.A(new_n634), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n465), .A2(G99gat), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n793), .B2(new_n811), .ZN(G1338gat));
  INV_X1    g611(.A(new_n785), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n710), .A2(new_n473), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(G106gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n473), .A2(new_n816), .A3(new_n634), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT114), .Z(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n791), .B2(new_n792), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n815), .A2(new_n821), .A3(new_n822), .A4(KEYINPUT53), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n816), .B1(new_n786), .B2(new_n473), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n820), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n823), .A2(new_n827), .ZN(G1339gat));
  NAND3_X1  g627(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(G229gat), .A3(G233gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n532), .B2(new_n535), .ZN(new_n831));
  INV_X1    g630(.A(new_n560), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n750), .A2(new_n634), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n608), .A2(new_n609), .A3(new_n613), .A4(new_n616), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n624), .B1(new_n836), .B2(new_n618), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n614), .A2(new_n629), .A3(new_n617), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n629), .B1(new_n614), .B2(new_n617), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n841), .A3(KEYINPUT55), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n837), .A2(new_n841), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n627), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT54), .B1(new_n628), .B2(new_n630), .ZN(new_n849));
  INV_X1    g648(.A(new_n618), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n623), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n848), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n844), .A2(new_n854), .A3(new_n627), .A4(new_n845), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n847), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n834), .B1(new_n856), .B2(new_n567), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n675), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n847), .A2(new_n855), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n750), .A2(new_n833), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n674), .A4(new_n853), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n661), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n660), .A2(new_n751), .A3(new_n634), .A4(new_n674), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n474), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n684), .A2(new_n430), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n567), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n567), .A2(G113gat), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT118), .Z(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n867), .B2(new_n870), .ZN(G1340gat));
  INV_X1    g670(.A(new_n867), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n634), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g673(.A1(new_n867), .A2(new_n660), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT119), .B(G127gat), .Z(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1342gat));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n674), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT56), .B(G134gat), .Z(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(G1343gat));
  OAI21_X1  g680(.A(new_n473), .B1(new_n862), .B2(new_n863), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n696), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n217), .B1(new_n886), .B2(new_n567), .ZN(new_n887));
  OR2_X1    g686(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n750), .A2(new_n634), .A3(new_n833), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n849), .B2(new_n852), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n837), .A2(new_n841), .A3(KEYINPUT120), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n848), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(new_n627), .A3(new_n844), .A4(new_n845), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n747), .B2(new_n750), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n675), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n861), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n863), .B1(new_n897), .B2(new_n660), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT57), .B1(new_n898), .B2(new_n259), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n473), .C1(new_n862), .C2(new_n863), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n567), .A2(new_n217), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n899), .A2(new_n901), .A3(new_n885), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n888), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n904), .B(new_n905), .ZN(G1344gat));
  NOR3_X1   g705(.A1(new_n469), .A2(new_n684), .A3(G148gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n883), .A2(new_n795), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n899), .A2(new_n901), .A3(new_n634), .A4(new_n885), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(G148gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n909), .A2(KEYINPUT122), .A3(new_n910), .A4(G148gat), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n863), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n896), .A2(new_n861), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n660), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n896), .B2(new_n861), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n900), .A3(new_n473), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n882), .A2(KEYINPUT57), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n922), .A2(new_n634), .A3(new_n885), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n910), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n908), .B1(new_n915), .B2(new_n925), .ZN(G1345gat));
  NAND3_X1  g725(.A1(new_n899), .A2(new_n885), .A3(new_n901), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n205), .A3(new_n660), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n886), .A2(new_n660), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n205), .ZN(G1346gat));
  NOR3_X1   g731(.A1(new_n927), .A2(new_n206), .A3(new_n675), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n883), .A2(new_n674), .A3(new_n885), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n206), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n428), .A2(new_n715), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n864), .A2(new_n474), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n567), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(new_n324), .ZN(G1348gat));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n810), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(new_n325), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n865), .A2(new_n352), .A3(new_n661), .A4(new_n936), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n314), .B(new_n315), .C1(new_n937), .C2(new_n660), .ZN(new_n943));
  NAND2_X1  g742(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g744(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(G1350gat));
  XNOR2_X1  g746(.A(KEYINPUT61), .B(G190gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n937), .A2(new_n675), .ZN(new_n950));
  MUX2_X1   g749(.A(new_n948), .B(new_n949), .S(new_n950), .Z(G1351gat));
  NAND2_X1  g750(.A1(new_n696), .A2(new_n936), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n922), .A2(new_n751), .A3(new_n923), .A4(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(G197gat), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n882), .A2(new_n952), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n751), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(G1352gat));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n620), .A3(new_n634), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n922), .A2(new_n923), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(new_n634), .A3(new_n953), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n964), .B(new_n965), .C1(new_n967), .C2(new_n620), .ZN(G1353gat));
  NAND4_X1  g767(.A1(new_n922), .A2(new_n661), .A3(new_n923), .A4(new_n953), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G211gat), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT63), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n959), .A2(new_n232), .A3(new_n661), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n971), .A2(KEYINPUT63), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(KEYINPUT63), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n969), .A2(G211gat), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(G1354gat));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n233), .A3(new_n674), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n966), .A2(new_n674), .A3(new_n953), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(new_n233), .ZN(G1355gat));
endmodule


