

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740;

  INV_X1 U375 ( .A(G146), .ZN(n428) );
  XNOR2_X1 U376 ( .A(n395), .B(KEYINPUT45), .ZN(n618) );
  XNOR2_X2 U377 ( .A(G122), .B(G113), .ZN(n410) );
  OR2_X2 U378 ( .A1(n622), .A2(G902), .ZN(n383) );
  XNOR2_X1 U379 ( .A(KEYINPUT85), .B(KEYINPUT3), .ZN(n411) );
  INV_X2 U380 ( .A(G953), .ZN(n732) );
  XNOR2_X1 U381 ( .A(n727), .B(n428), .ZN(n367) );
  NOR2_X1 U382 ( .A1(n740), .A2(n739), .ZN(n415) );
  XNOR2_X1 U383 ( .A(n603), .B(n602), .ZN(n739) );
  OR2_X1 U384 ( .A1(n611), .A2(n673), .ZN(n603) );
  XNOR2_X1 U385 ( .A(n375), .B(KEYINPUT39), .ZN(n611) );
  AND2_X1 U386 ( .A1(n374), .A2(n574), .ZN(n375) );
  AND2_X1 U387 ( .A1(n527), .A2(n526), .ZN(n557) );
  XNOR2_X1 U388 ( .A(KEYINPUT62), .B(n632), .ZN(n421) );
  XNOR2_X1 U389 ( .A(n483), .B(n367), .ZN(n632) );
  XNOR2_X1 U390 ( .A(n435), .B(n427), .ZN(n727) );
  XNOR2_X1 U391 ( .A(n410), .B(n441), .ZN(n382) );
  XNOR2_X1 U392 ( .A(n499), .B(G134), .ZN(n435) );
  NOR2_X1 U393 ( .A1(n621), .A2(n687), .ZN(n353) );
  NOR2_X2 U394 ( .A1(n621), .A2(n687), .ZN(n354) );
  BUF_X1 U395 ( .A(n585), .Z(n355) );
  NOR2_X2 U396 ( .A1(n621), .A2(n687), .ZN(n646) );
  NOR2_X4 U397 ( .A1(n620), .A2(n619), .ZN(n687) );
  BUF_X1 U398 ( .A(n599), .Z(n576) );
  XNOR2_X2 U399 ( .A(G143), .B(G128), .ZN(n499) );
  XNOR2_X1 U400 ( .A(n605), .B(n390), .ZN(n708) );
  INV_X1 U401 ( .A(KEYINPUT111), .ZN(n390) );
  XNOR2_X1 U402 ( .A(n465), .B(n464), .ZN(n527) );
  XNOR2_X1 U403 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U404 ( .A(n518), .B(n517), .ZN(n521) );
  XNOR2_X1 U405 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n517) );
  XNOR2_X1 U406 ( .A(n497), .B(n443), .ZN(n455) );
  XNOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n443) );
  XNOR2_X1 U408 ( .A(n495), .B(n496), .ZN(n386) );
  XNOR2_X1 U409 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n496) );
  XNOR2_X1 U410 ( .A(n428), .B(G125), .ZN(n497) );
  XNOR2_X1 U411 ( .A(n369), .B(n391), .ZN(n368) );
  INV_X1 U412 ( .A(KEYINPUT48), .ZN(n391) );
  AND2_X1 U413 ( .A1(n610), .A2(n356), .ZN(n416) );
  XNOR2_X1 U414 ( .A(n440), .B(n439), .ZN(n534) );
  NOR2_X1 U415 ( .A1(G902), .A2(n650), .ZN(n440) );
  XNOR2_X1 U416 ( .A(G116), .B(G107), .ZN(n494) );
  XNOR2_X1 U417 ( .A(n457), .B(n401), .ZN(n400) );
  XNOR2_X1 U418 ( .A(G119), .B(G128), .ZN(n457) );
  XNOR2_X1 U419 ( .A(n402), .B(KEYINPUT89), .ZN(n401) );
  INV_X1 U420 ( .A(KEYINPUT24), .ZN(n402) );
  XNOR2_X1 U421 ( .A(n432), .B(n419), .ZN(n456) );
  INV_X1 U422 ( .A(KEYINPUT8), .ZN(n419) );
  XNOR2_X1 U423 ( .A(n455), .B(n454), .ZN(n726) );
  NAND2_X1 U424 ( .A1(n456), .A2(G217), .ZN(n418) );
  XNOR2_X1 U425 ( .A(n494), .B(G122), .ZN(n417) );
  NOR2_X1 U426 ( .A1(n708), .A2(n604), .ZN(n607) );
  XNOR2_X1 U427 ( .A(n429), .B(G469), .ZN(n430) );
  INV_X1 U428 ( .A(n658), .ZN(n634) );
  NOR2_X1 U429 ( .A1(n725), .A2(n724), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n407), .B(n406), .ZN(n543) );
  INV_X1 U431 ( .A(KEYINPUT107), .ZN(n406) );
  INV_X1 U432 ( .A(KEYINPUT69), .ZN(n547) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n466) );
  INV_X1 U434 ( .A(G237), .ZN(n490) );
  XNOR2_X1 U435 ( .A(n405), .B(n530), .ZN(n531) );
  NOR2_X1 U436 ( .A1(n397), .A2(n525), .ZN(n405) );
  INV_X1 U437 ( .A(n557), .ZN(n693) );
  XNOR2_X1 U438 ( .A(G137), .B(G116), .ZN(n478) );
  XOR2_X1 U439 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n477) );
  AND2_X1 U440 ( .A1(n368), .A2(n613), .ZN(n730) );
  XNOR2_X1 U441 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n409) );
  INV_X1 U442 ( .A(G104), .ZN(n441) );
  XNOR2_X1 U443 ( .A(n412), .B(n411), .ZN(n381) );
  XNOR2_X1 U444 ( .A(G119), .B(G101), .ZN(n412) );
  XNOR2_X1 U445 ( .A(G101), .B(G107), .ZN(n422) );
  XOR2_X1 U446 ( .A(G110), .B(G104), .Z(n423) );
  XNOR2_X1 U447 ( .A(n384), .B(n500), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n497), .ZN(n384) );
  NAND2_X1 U449 ( .A1(n368), .A2(n359), .ZN(n617) );
  XNOR2_X1 U450 ( .A(n378), .B(n377), .ZN(n585) );
  INV_X1 U451 ( .A(KEYINPUT19), .ZN(n377) );
  XNOR2_X1 U452 ( .A(n413), .B(KEYINPUT30), .ZN(n574) );
  NOR2_X1 U453 ( .A1(n582), .A2(n508), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n519), .B(KEYINPUT106), .ZN(n582) );
  XNOR2_X1 U455 ( .A(n389), .B(n387), .ZN(n408) );
  XNOR2_X1 U456 ( .A(n388), .B(n494), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n381), .B(n382), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n409), .B(G110), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n398), .B(n726), .ZN(n648) );
  XNOR2_X1 U460 ( .A(n459), .B(n399), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n458), .B(n400), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n438), .B(n437), .ZN(n650) );
  XNOR2_X1 U463 ( .A(n418), .B(n417), .ZN(n438) );
  XNOR2_X1 U464 ( .A(KEYINPUT42), .B(n609), .ZN(n740) );
  NAND2_X1 U465 ( .A1(n404), .A2(n420), .ZN(n403) );
  INV_X1 U466 ( .A(KEYINPUT56), .ZN(n392) );
  XNOR2_X1 U467 ( .A(n371), .B(n370), .ZN(G75) );
  INV_X1 U468 ( .A(KEYINPUT53), .ZN(n370) );
  XNOR2_X1 U469 ( .A(n373), .B(KEYINPUT122), .ZN(n372) );
  INV_X1 U470 ( .A(n543), .ZN(n542) );
  AND2_X1 U471 ( .A1(n669), .A2(n587), .ZN(n356) );
  XOR2_X1 U472 ( .A(n426), .B(n425), .Z(n357) );
  XOR2_X1 U473 ( .A(n453), .B(G475), .Z(n358) );
  AND2_X1 U474 ( .A1(n613), .A2(KEYINPUT2), .ZN(n359) );
  AND2_X1 U475 ( .A1(n600), .A2(n705), .ZN(n360) );
  AND2_X1 U476 ( .A1(n582), .A2(n520), .ZN(n361) );
  NOR2_X1 U477 ( .A1(n588), .A2(n380), .ZN(n362) );
  XOR2_X1 U478 ( .A(n379), .B(n628), .Z(n363) );
  XNOR2_X1 U479 ( .A(KEYINPUT59), .B(n622), .ZN(n364) );
  NOR2_X1 U480 ( .A1(n408), .A2(n644), .ZN(n365) );
  XNOR2_X1 U481 ( .A(n625), .B(KEYINPUT65), .ZN(n366) );
  XNOR2_X1 U482 ( .A(n357), .B(n367), .ZN(n655) );
  NAND2_X1 U483 ( .A1(n414), .A2(n416), .ZN(n369) );
  NAND2_X1 U484 ( .A1(n372), .A2(n732), .ZN(n371) );
  NAND2_X1 U485 ( .A1(n574), .A2(n575), .ZN(n601) );
  AND2_X1 U486 ( .A1(n575), .A2(n360), .ZN(n374) );
  XNOR2_X2 U487 ( .A(n376), .B(n515), .ZN(n553) );
  NAND2_X1 U488 ( .A1(n585), .A2(n513), .ZN(n376) );
  NOR2_X2 U489 ( .A1(n599), .A2(n508), .ZN(n378) );
  BUF_X1 U490 ( .A(n629), .Z(n379) );
  OR2_X1 U491 ( .A1(n576), .A2(n508), .ZN(n380) );
  XNOR2_X1 U492 ( .A(n381), .B(n482), .ZN(n483) );
  XNOR2_X1 U493 ( .A(n382), .B(n442), .ZN(n444) );
  XNOR2_X1 U494 ( .A(n452), .B(n451), .ZN(n622) );
  NOR2_X1 U495 ( .A1(n562), .A2(n534), .ZN(n506) );
  XNOR2_X2 U496 ( .A(n383), .B(n358), .ZN(n562) );
  XNOR2_X1 U497 ( .A(n408), .B(n385), .ZN(n629) );
  NAND2_X1 U498 ( .A1(n556), .A2(n531), .ZN(n533) );
  XNOR2_X1 U499 ( .A(n393), .B(n392), .ZN(G51) );
  NAND2_X1 U500 ( .A1(n631), .A2(n634), .ZN(n393) );
  XNOR2_X1 U501 ( .A(n394), .B(n366), .ZN(G60) );
  NAND2_X1 U502 ( .A1(n624), .A2(n634), .ZN(n394) );
  NAND2_X1 U503 ( .A1(n571), .A2(n572), .ZN(n395) );
  XNOR2_X1 U504 ( .A(n396), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U505 ( .A1(n635), .A2(n634), .ZN(n396) );
  XNOR2_X2 U506 ( .A(n504), .B(n503), .ZN(n599) );
  XNOR2_X1 U507 ( .A(n600), .B(KEYINPUT1), .ZN(n528) );
  XNOR2_X2 U508 ( .A(n431), .B(n430), .ZN(n600) );
  NAND2_X1 U509 ( .A1(n528), .A2(n557), .ZN(n397) );
  NAND2_X1 U510 ( .A1(n544), .A2(n543), .ZN(n549) );
  XNOR2_X2 U511 ( .A(n403), .B(KEYINPUT32), .ZN(n544) );
  INV_X1 U512 ( .A(n541), .ZN(n404) );
  INV_X1 U513 ( .A(n525), .ZN(n488) );
  INV_X1 U514 ( .A(n531), .ZN(n719) );
  INV_X1 U515 ( .A(n544), .ZN(n637) );
  NAND2_X1 U516 ( .A1(n521), .A2(n361), .ZN(n407) );
  NAND2_X1 U517 ( .A1(n553), .A2(n516), .ZN(n518) );
  XNOR2_X1 U518 ( .A(n553), .B(KEYINPUT88), .ZN(n556) );
  XNOR2_X1 U519 ( .A(n415), .B(KEYINPUT46), .ZN(n414) );
  BUF_X1 U520 ( .A(n618), .Z(n639) );
  AND2_X1 U521 ( .A1(n688), .A2(n589), .ZN(n420) );
  NOR2_X1 U522 ( .A1(n732), .A2(G952), .ZN(n658) );
  XNOR2_X1 U523 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U524 ( .A(G131), .B(KEYINPUT4), .ZN(n427) );
  INV_X1 U525 ( .A(G478), .ZN(n439) );
  XNOR2_X1 U526 ( .A(G137), .B(G140), .ZN(n454) );
  XNOR2_X1 U527 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U528 ( .A(n454), .B(n424), .ZN(n426) );
  NAND2_X1 U529 ( .A1(G227), .A2(n732), .ZN(n425) );
  NOR2_X1 U530 ( .A1(n655), .A2(G902), .ZN(n431) );
  INV_X1 U531 ( .A(KEYINPUT68), .ZN(n429) );
  BUF_X1 U532 ( .A(n528), .Z(n589) );
  NAND2_X1 U533 ( .A1(G234), .A2(n732), .ZN(n432) );
  XOR2_X1 U534 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n434) );
  XNOR2_X1 U535 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n433) );
  XNOR2_X1 U536 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U537 ( .A(n435), .B(n436), .ZN(n437) );
  INV_X1 U538 ( .A(n534), .ZN(n561) );
  NOR2_X1 U539 ( .A1(G953), .A2(G237), .ZN(n475) );
  NAND2_X1 U540 ( .A1(G214), .A2(n475), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n444), .B(n455), .ZN(n452) );
  XOR2_X1 U542 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n446) );
  XNOR2_X1 U543 ( .A(G143), .B(G131), .ZN(n445) );
  XNOR2_X1 U544 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U545 ( .A(G140), .B(KEYINPUT12), .Z(n448) );
  XNOR2_X1 U546 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n447) );
  XNOR2_X1 U547 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U548 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U549 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n453) );
  NAND2_X1 U550 ( .A1(n561), .A2(n562), .ZN(n673) );
  AND2_X1 U551 ( .A1(n456), .A2(G221), .ZN(n459) );
  XOR2_X1 U552 ( .A(KEYINPUT23), .B(G110), .Z(n458) );
  NOR2_X1 U553 ( .A1(G902), .A2(n648), .ZN(n465) );
  XNOR2_X1 U554 ( .A(G902), .B(KEYINPUT15), .ZN(n501) );
  NAND2_X1 U555 ( .A1(G234), .A2(n501), .ZN(n460) );
  XNOR2_X1 U556 ( .A(KEYINPUT20), .B(n460), .ZN(n472) );
  AND2_X1 U557 ( .A1(n472), .A2(G217), .ZN(n461) );
  XNOR2_X1 U558 ( .A(n461), .B(KEYINPUT91), .ZN(n463) );
  XNOR2_X1 U559 ( .A(KEYINPUT25), .B(KEYINPUT90), .ZN(n462) );
  XNOR2_X1 U560 ( .A(n466), .B(KEYINPUT86), .ZN(n467) );
  XNOR2_X1 U561 ( .A(KEYINPUT14), .B(n467), .ZN(n468) );
  NAND2_X1 U562 ( .A1(G952), .A2(n468), .ZN(n717) );
  NOR2_X1 U563 ( .A1(n717), .A2(G953), .ZN(n511) );
  AND2_X1 U564 ( .A1(n468), .A2(G902), .ZN(n509) );
  NAND2_X1 U565 ( .A1(G953), .A2(n509), .ZN(n469) );
  NOR2_X1 U566 ( .A1(G900), .A2(n469), .ZN(n470) );
  NOR2_X1 U567 ( .A1(n511), .A2(n470), .ZN(n471) );
  XOR2_X1 U568 ( .A(KEYINPUT75), .B(n471), .Z(n573) );
  NOR2_X1 U569 ( .A1(n527), .A2(n573), .ZN(n474) );
  NAND2_X1 U570 ( .A1(n472), .A2(G221), .ZN(n473) );
  XNOR2_X1 U571 ( .A(n473), .B(KEYINPUT21), .ZN(n689) );
  INV_X1 U572 ( .A(n689), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n474), .A2(n526), .ZN(n581) );
  NOR2_X1 U574 ( .A1(n673), .A2(n581), .ZN(n489) );
  NAND2_X1 U575 ( .A1(n475), .A2(G210), .ZN(n476) );
  XNOR2_X1 U576 ( .A(n477), .B(n476), .ZN(n481) );
  XOR2_X1 U577 ( .A(KEYINPUT93), .B(G113), .Z(n479) );
  XNOR2_X1 U578 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U579 ( .A(G902), .ZN(n491) );
  NAND2_X1 U580 ( .A1(n632), .A2(n491), .ZN(n485) );
  XOR2_X1 U581 ( .A(G472), .B(KEYINPUT70), .Z(n484) );
  XNOR2_X2 U582 ( .A(n485), .B(n484), .ZN(n519) );
  INV_X1 U583 ( .A(n519), .ZN(n558) );
  INV_X1 U584 ( .A(KEYINPUT102), .ZN(n486) );
  XNOR2_X1 U585 ( .A(n486), .B(KEYINPUT6), .ZN(n487) );
  XNOR2_X1 U586 ( .A(n519), .B(n487), .ZN(n525) );
  NAND2_X1 U587 ( .A1(n489), .A2(n488), .ZN(n588) );
  NOR2_X1 U588 ( .A1(n589), .A2(n588), .ZN(n492) );
  NAND2_X1 U589 ( .A1(n491), .A2(n490), .ZN(n502) );
  NAND2_X1 U590 ( .A1(n502), .A2(G214), .ZN(n704) );
  NAND2_X1 U591 ( .A1(n492), .A2(n704), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n493), .B(KEYINPUT43), .ZN(n505) );
  NAND2_X1 U593 ( .A1(n732), .A2(G224), .ZN(n495) );
  XNOR2_X1 U594 ( .A(KEYINPUT73), .B(KEYINPUT4), .ZN(n498) );
  XNOR2_X1 U595 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U596 ( .A(n501), .ZN(n614) );
  OR2_X2 U597 ( .A1(n629), .A2(n614), .ZN(n504) );
  NAND2_X1 U598 ( .A1(n502), .A2(G210), .ZN(n503) );
  AND2_X1 U599 ( .A1(n505), .A2(n576), .ZN(n612) );
  XOR2_X1 U600 ( .A(n612), .B(G140), .Z(G42) );
  XNOR2_X1 U601 ( .A(n506), .B(KEYINPUT103), .ZN(n604) );
  NOR2_X1 U602 ( .A1(n604), .A2(n689), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n507), .B(KEYINPUT104), .ZN(n516) );
  INV_X1 U604 ( .A(n704), .ZN(n508) );
  NOR2_X1 U605 ( .A1(G898), .A2(n732), .ZN(n644) );
  NAND2_X1 U606 ( .A1(n644), .A2(n509), .ZN(n510) );
  XNOR2_X1 U607 ( .A(n510), .B(KEYINPUT87), .ZN(n512) );
  OR2_X1 U608 ( .A1(n512), .A2(n511), .ZN(n513) );
  INV_X1 U609 ( .A(KEYINPUT84), .ZN(n514) );
  XNOR2_X1 U610 ( .A(n514), .B(KEYINPUT0), .ZN(n515) );
  NOR2_X1 U611 ( .A1(n589), .A2(n527), .ZN(n520) );
  XOR2_X1 U612 ( .A(G110), .B(n542), .Z(G12) );
  NAND2_X1 U613 ( .A1(n521), .A2(n525), .ZN(n541) );
  NOR2_X1 U614 ( .A1(n541), .A2(n589), .ZN(n522) );
  XOR2_X1 U615 ( .A(KEYINPUT79), .B(n522), .Z(n524) );
  XNOR2_X1 U616 ( .A(n527), .B(KEYINPUT105), .ZN(n688) );
  INV_X1 U617 ( .A(n688), .ZN(n523) );
  NAND2_X1 U618 ( .A1(n524), .A2(n523), .ZN(n567) );
  XNOR2_X1 U619 ( .A(n567), .B(G101), .ZN(G3) );
  INV_X1 U620 ( .A(KEYINPUT108), .ZN(n529) );
  XNOR2_X1 U621 ( .A(n529), .B(KEYINPUT33), .ZN(n530) );
  INV_X1 U622 ( .A(KEYINPUT34), .ZN(n532) );
  XNOR2_X1 U623 ( .A(n533), .B(n532), .ZN(n537) );
  AND2_X1 U624 ( .A1(n562), .A2(n534), .ZN(n536) );
  INV_X1 U625 ( .A(KEYINPUT109), .ZN(n535) );
  XNOR2_X1 U626 ( .A(n536), .B(n535), .ZN(n580) );
  NAND2_X1 U627 ( .A1(n537), .A2(n580), .ZN(n539) );
  XNOR2_X1 U628 ( .A(KEYINPUT74), .B(KEYINPUT35), .ZN(n538) );
  XNOR2_X2 U629 ( .A(n539), .B(n538), .ZN(n638) );
  NOR2_X2 U630 ( .A1(n638), .A2(KEYINPUT44), .ZN(n540) );
  XNOR2_X1 U631 ( .A(n540), .B(KEYINPUT66), .ZN(n546) );
  XNOR2_X1 U632 ( .A(n549), .B(KEYINPUT81), .ZN(n545) );
  NAND2_X1 U633 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U634 ( .A(n548), .B(n547), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n549), .A2(n638), .ZN(n551) );
  INV_X1 U636 ( .A(KEYINPUT44), .ZN(n550) );
  NOR2_X1 U637 ( .A1(n551), .A2(n550), .ZN(n569) );
  INV_X1 U638 ( .A(n589), .ZN(n692) );
  NAND2_X1 U639 ( .A1(n558), .A2(n557), .ZN(n552) );
  NOR2_X1 U640 ( .A1(n692), .A2(n552), .ZN(n701) );
  NAND2_X1 U641 ( .A1(n701), .A2(n553), .ZN(n555) );
  XOR2_X1 U642 ( .A(KEYINPUT31), .B(KEYINPUT94), .Z(n554) );
  XNOR2_X1 U643 ( .A(n555), .B(n554), .ZN(n677) );
  NAND2_X1 U644 ( .A1(n557), .A2(n600), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n556), .A2(n560), .ZN(n662) );
  NAND2_X1 U647 ( .A1(n677), .A2(n662), .ZN(n565) );
  NOR2_X1 U648 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U649 ( .A(n563), .B(KEYINPUT101), .ZN(n676) );
  NAND2_X1 U650 ( .A1(n673), .A2(n676), .ZN(n707) );
  XNOR2_X1 U651 ( .A(KEYINPUT76), .B(n707), .ZN(n564) );
  NAND2_X1 U652 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U653 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X2 U654 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U655 ( .A(n570), .B(KEYINPUT80), .ZN(n571) );
  NOR2_X1 U656 ( .A1(n573), .A2(n693), .ZN(n575) );
  INV_X1 U657 ( .A(n576), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n600), .A2(n577), .ZN(n578) );
  NOR2_X1 U659 ( .A1(n601), .A2(n578), .ZN(n579) );
  NAND2_X1 U660 ( .A1(n580), .A2(n579), .ZN(n669) );
  NOR2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U662 ( .A(KEYINPUT28), .B(n583), .ZN(n584) );
  NAND2_X1 U663 ( .A1(n584), .A2(n600), .ZN(n608) );
  INV_X1 U664 ( .A(n355), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n608), .A2(n586), .ZN(n671) );
  INV_X1 U666 ( .A(n671), .ZN(n666) );
  NAND2_X1 U667 ( .A1(n666), .A2(KEYINPUT47), .ZN(n587) );
  XNOR2_X1 U668 ( .A(n362), .B(KEYINPUT36), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n681) );
  XNOR2_X1 U670 ( .A(KEYINPUT78), .B(n681), .ZN(n594) );
  NAND2_X1 U671 ( .A1(KEYINPUT76), .A2(n707), .ZN(n591) );
  NOR2_X1 U672 ( .A1(n591), .A2(KEYINPUT47), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n671), .A2(n592), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n598) );
  NOR2_X1 U675 ( .A1(n666), .A2(KEYINPUT76), .ZN(n595) );
  NOR2_X1 U676 ( .A1(KEYINPUT47), .A2(n595), .ZN(n596) );
  NOR2_X1 U677 ( .A1(n596), .A2(n707), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n598), .A2(n597), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n576), .B(KEYINPUT38), .ZN(n705) );
  XOR2_X1 U680 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n602) );
  NAND2_X1 U681 ( .A1(n705), .A2(n704), .ZN(n605) );
  XNOR2_X1 U682 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n607), .B(n606), .ZN(n718) );
  NOR2_X1 U684 ( .A1(n718), .A2(n608), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n611), .A2(n676), .ZN(n683) );
  NOR2_X1 U686 ( .A1(n683), .A2(n612), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n618), .A2(n730), .ZN(n685) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n684) );
  NAND2_X1 U689 ( .A1(n685), .A2(n684), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X2 U691 ( .A(n616), .B(KEYINPUT64), .ZN(n621) );
  XOR2_X1 U692 ( .A(n617), .B(KEYINPUT77), .Z(n620) );
  INV_X1 U693 ( .A(n639), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n646), .A2(G475), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(n364), .ZN(n624) );
  XNOR2_X1 U696 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n646), .A2(G210), .ZN(n630) );
  XNOR2_X1 U698 ( .A(KEYINPUT83), .B(KEYINPUT54), .ZN(n627) );
  XNOR2_X1 U699 ( .A(KEYINPUT55), .B(KEYINPUT82), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n630), .B(n363), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n354), .A2(G472), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(n421), .ZN(n635) );
  XNOR2_X1 U704 ( .A(G119), .B(KEYINPUT127), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(G21) );
  XOR2_X1 U706 ( .A(n638), .B(G122), .Z(G24) );
  NAND2_X1 U707 ( .A1(n639), .A2(n732), .ZN(n643) );
  NAND2_X1 U708 ( .A1(G953), .A2(G224), .ZN(n640) );
  XNOR2_X1 U709 ( .A(KEYINPUT61), .B(n640), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n641), .A2(G898), .ZN(n642) );
  NAND2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n645) );
  XNOR2_X1 U712 ( .A(n645), .B(n365), .ZN(G69) );
  NAND2_X1 U713 ( .A1(n353), .A2(G217), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U715 ( .A1(n649), .A2(n658), .ZN(G66) );
  NAND2_X1 U716 ( .A1(n354), .A2(G478), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n652), .A2(n658), .ZN(G63) );
  NAND2_X1 U719 ( .A1(n353), .A2(G469), .ZN(n657) );
  XNOR2_X1 U720 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT58), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U723 ( .A(n657), .B(n656), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(G54) );
  NOR2_X1 U725 ( .A1(n662), .A2(n673), .ZN(n661) );
  XNOR2_X1 U726 ( .A(G104), .B(KEYINPUT113), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n661), .B(n660), .ZN(G6) );
  NOR2_X1 U728 ( .A1(n662), .A2(n676), .ZN(n664) );
  XNOR2_X1 U729 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U731 ( .A(G107), .B(n665), .ZN(G9) );
  NOR2_X1 U732 ( .A1(n666), .A2(n676), .ZN(n668) );
  XNOR2_X1 U733 ( .A(G128), .B(KEYINPUT29), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n668), .B(n667), .ZN(G30) );
  XNOR2_X1 U735 ( .A(G143), .B(n669), .ZN(G45) );
  INV_X1 U736 ( .A(n673), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(G146), .ZN(G48) );
  NOR2_X1 U739 ( .A1(n677), .A2(n673), .ZN(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT114), .B(n674), .Z(n675) );
  XNOR2_X1 U741 ( .A(G113), .B(n675), .ZN(G15) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U743 ( .A(G116), .B(KEYINPUT115), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n679), .B(n678), .ZN(G18) );
  XOR2_X1 U745 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n680) );
  XNOR2_X1 U746 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U747 ( .A(G125), .B(n682), .ZN(G27) );
  XOR2_X1 U748 ( .A(G134), .B(n683), .Z(G36) );
  AND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n725) );
  XOR2_X1 U751 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n691) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n691), .B(n690), .ZN(n699) );
  XOR2_X1 U754 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n695) );
  NAND2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(KEYINPUT118), .B(n696), .ZN(n697) );
  NAND2_X1 U758 ( .A1(n697), .A2(n519), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U761 ( .A(KEYINPUT51), .B(n702), .Z(n703) );
  NOR2_X1 U762 ( .A1(n718), .A2(n703), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n604), .A2(n706), .ZN(n711) );
  INV_X1 U765 ( .A(n707), .ZN(n709) );
  NOR2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U768 ( .A1(n719), .A2(n712), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U770 ( .A(n715), .B(KEYINPUT52), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n722) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT120), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n723), .B(KEYINPUT121), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n728), .B(KEYINPUT125), .ZN(n734) );
  INV_X1 U778 ( .A(n734), .ZN(n729) );
  XNOR2_X1 U779 ( .A(KEYINPUT126), .B(n729), .ZN(n731) );
  XNOR2_X1 U780 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(n738) );
  XNOR2_X1 U782 ( .A(G227), .B(n734), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(G900), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G953), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n738), .A2(n737), .ZN(G72) );
  XOR2_X1 U786 ( .A(n739), .B(G131), .Z(G33) );
  XOR2_X1 U787 ( .A(n740), .B(G137), .Z(G39) );
endmodule

