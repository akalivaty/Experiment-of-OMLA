//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT66), .B(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n467), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(G124), .A2(new_n477), .B1(new_n478), .B2(G136), .ZN(new_n479));
  OAI221_X1 g054(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n484), .B(new_n485), .C1(new_n472), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n465), .A2(G102), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n487), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n484), .B1(new_n472), .B2(new_n486), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n460), .A3(KEYINPUT68), .A4(G138), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n483), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n490), .A2(G2105), .B1(G102), .B2(new_n465), .ZN(new_n498));
  AND4_X1   g073(.A1(new_n483), .A2(new_n496), .A3(new_n487), .A4(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n509), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT70), .ZN(new_n519));
  INV_X1    g094(.A(new_n514), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(new_n511), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n519), .A2(new_n521), .A3(new_n523), .A4(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n508), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n511), .A2(new_n530), .B1(new_n531), .B2(new_n514), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G171));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n503), .A2(new_n505), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT71), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(new_n541), .B1(G43), .B2(new_n520), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT73), .B(G81), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n524), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n520), .A2(G53), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n553), .B(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G91), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n508), .B1(new_n511), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n556), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  NAND2_X1  g136(.A1(new_n524), .A2(G87), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n520), .A2(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND3_X1  g140(.A1(new_n506), .A2(KEYINPUT75), .A3(G61), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n535), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G48), .B2(new_n520), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n524), .A2(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G305));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n511), .A2(new_n575), .B1(new_n576), .B2(new_n514), .ZN(new_n577));
  NAND2_X1  g152(.A1(G72), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G60), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n535), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n577), .B1(G651), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  INV_X1    g158(.A(G92), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n511), .A2(KEYINPUT10), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT10), .B1(new_n511), .B2(new_n584), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n508), .B1(new_n514), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n583), .B1(G868), .B2(new_n591), .ZN(G284));
  OAI21_X1  g167(.A(new_n583), .B1(G868), .B2(new_n591), .ZN(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n556), .A2(new_n559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n591), .B1(new_n598), .B2(G860), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT77), .Z(G148));
  INV_X1    g175(.A(new_n591), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(G559), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n546), .B2(G868), .ZN(G323));
  XOR2_X1   g180(.A(G323), .B(KEYINPUT78), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n477), .A2(G123), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n478), .A2(G135), .ZN(new_n609));
  OAI221_X1 g184(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  XOR2_X1   g187(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n613));
  NOR3_X1   g188(.A1(new_n468), .A2(new_n464), .A3(G2105), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G2100), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n615), .B(new_n618), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n612), .B(new_n619), .C1(new_n616), .C2(G2100), .ZN(G156));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2427), .B(G2430), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n632), .B(new_n633), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G14), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n637), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  AOI21_X1  g221(.A(KEYINPUT18), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n644), .B(new_n647), .Z(G227));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XOR2_X1   g226(.A(G1961), .B(G1966), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT83), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT20), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n650), .A3(new_n653), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n659), .C1(new_n650), .C2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT22), .B(G1981), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G229));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n668));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n669), .A2(G6), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(G305), .B2(G16), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT32), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT86), .B(G1981), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n669), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n669), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(KEYINPUT33), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(KEYINPUT33), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G1976), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n669), .A2(G22), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n669), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G1971), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(G1976), .A3(new_n682), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n687), .A2(G1971), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n677), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n668), .B1(new_n692), .B2(KEYINPUT34), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n690), .A2(new_n677), .A3(new_n694), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n477), .A2(G119), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT84), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n478), .A2(G131), .ZN(new_n698));
  OAI221_X1 g273(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G25), .B(new_n700), .S(G29), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT35), .B(G1991), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  MUX2_X1   g278(.A(G24), .B(G290), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT85), .B(G1986), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n693), .A2(new_n695), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n669), .A2(KEYINPUT23), .A3(G20), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT23), .ZN(new_n711));
  INV_X1    g286(.A(G20), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n713), .C1(new_n595), .C2(new_n669), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1956), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  AOI22_X1  g292(.A1(G129), .A2(new_n477), .B1(new_n478), .B2(G141), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n465), .A2(G105), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT26), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G32), .B(new_n724), .S(G29), .Z(new_n725));
  AOI21_X1  g300(.A(new_n715), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n727), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n731));
  OAI21_X1  g306(.A(G2090), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n733));
  INV_X1    g308(.A(new_n478), .ZN(new_n734));
  INV_X1    g309(.A(G140), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n477), .A2(G128), .ZN(new_n737));
  OAI221_X1 g312(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n478), .A2(KEYINPUT88), .A3(G140), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n727), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT90), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2067), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n727), .B1(new_n748), .B2(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(G28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AND4_X1   g328(.A1(new_n726), .A2(new_n732), .A3(new_n747), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n727), .A2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G139), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n758), .B1(new_n759), .B2(new_n734), .C1(new_n462), .C2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n755), .B1(new_n762), .B2(new_n727), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G2072), .Z(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT31), .B(G11), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n669), .A2(G5), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G171), .B2(new_n669), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1961), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n669), .A2(G21), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G286), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(KEYINPUT24), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(KEYINPUT24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n727), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n727), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2084), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n591), .B2(G16), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n779), .B1(new_n771), .B2(new_n772), .C1(new_n781), .C2(G1348), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n766), .A2(new_n769), .A3(new_n773), .A4(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n725), .A2(new_n717), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n781), .A2(G1348), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n669), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n545), .B2(G16), .ZN(new_n791));
  INV_X1    g366(.A(G1341), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n730), .A2(new_n731), .A3(G2090), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n754), .A2(new_n783), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n707), .B2(new_n708), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n611), .A2(new_n727), .ZN(new_n799));
  NOR2_X1   g374(.A1(G27), .A2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(G29), .ZN(new_n801));
  INV_X1    g376(.A(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n709), .A2(new_n798), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n778), .A2(G2084), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(G311));
  AND3_X1   g381(.A1(new_n709), .A2(new_n803), .A3(new_n798), .ZN(new_n807));
  INV_X1    g382(.A(new_n805), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n807), .A2(KEYINPUT96), .A3(new_n808), .A4(new_n799), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n804), .B2(new_n805), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(G150));
  AOI22_X1  g387(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n508), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n511), .A2(new_n815), .B1(new_n816), .B2(new_n514), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n546), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n545), .A2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n601), .A2(new_n598), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT97), .ZN(new_n828));
  AOI21_X1  g403(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(KEYINPUT97), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n819), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(G145));
  AOI22_X1  g409(.A1(G130), .A2(new_n477), .B1(new_n478), .B2(G142), .ZN(new_n835));
  OAI221_X1 g410(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n462), .C2(G118), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n615), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n700), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n496), .A2(new_n487), .A3(new_n498), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n740), .B(new_n841), .Z(new_n842));
  OR2_X1    g417(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n761), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n762), .A2(new_n722), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n845), .A2(new_n842), .A3(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(new_n839), .A3(new_n847), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT99), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(G160), .B(new_n611), .Z(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(G162), .Z(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n850), .B2(KEYINPUT99), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n852), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n839), .B1(new_n851), .B2(new_n847), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(KEYINPUT100), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  INV_X1    g438(.A(new_n856), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n861), .B(new_n863), .C1(new_n853), .C2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g446(.A1(new_n819), .A2(G868), .ZN(new_n872));
  NAND2_X1  g447(.A1(G299), .A2(new_n591), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n601), .A2(new_n595), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n601), .B2(new_n595), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n875), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n877), .B1(new_n880), .B2(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n820), .B2(new_n821), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n820), .A2(new_n883), .A3(new_n821), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n602), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n602), .A3(new_n886), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n891), .A2(new_n887), .A3(new_n876), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT106), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(G288), .B(KEYINPUT103), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G290), .ZN(new_n895));
  XNOR2_X1  g470(.A(G305), .B(G303), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(KEYINPUT105), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n881), .B1(new_n891), .B2(new_n887), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n888), .A2(new_n889), .A3(new_n875), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n905), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n893), .A2(new_n907), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n890), .A2(new_n892), .ZN(new_n914));
  INV_X1    g489(.A(new_n912), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n914), .B(new_n910), .C1(new_n915), .C2(new_n906), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n872), .B1(new_n917), .B2(G868), .ZN(G295));
  AOI21_X1  g493(.A(new_n872), .B1(new_n917), .B2(G868), .ZN(G331));
  XNOR2_X1  g494(.A(G286), .B(G301), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n822), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n820), .A2(new_n821), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n881), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n875), .A3(new_n923), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n903), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n863), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n875), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n880), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n903), .B1(new_n937), .B2(new_n926), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n928), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n903), .B1(new_n925), .B2(new_n926), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n928), .A2(KEYINPUT43), .A3(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(KEYINPUT109), .B(KEYINPUT43), .C1(new_n928), .C2(new_n938), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n941), .A2(KEYINPUT44), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n928), .B2(new_n942), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n928), .A2(KEYINPUT43), .A3(new_n938), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(KEYINPUT44), .B2(new_n949), .ZN(G397));
  AOI21_X1  g525(.A(G1384), .B1(new_n493), .B2(new_n496), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(KEYINPUT45), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G160), .A2(G40), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n953), .A2(KEYINPUT110), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OR3_X1    g532(.A1(new_n957), .A2(G1986), .A3(G290), .ZN(new_n958));
  INV_X1    g533(.A(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G1986), .A3(G290), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT111), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n740), .B(G2067), .Z(new_n963));
  NAND2_X1  g538(.A1(new_n722), .A2(G1996), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n963), .B(new_n964), .C1(new_n724), .C2(G1996), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n700), .A2(new_n702), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n700), .A2(new_n702), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n959), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n962), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT121), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n559), .B2(KEYINPUT120), .ZN(new_n973));
  XNOR2_X1  g548(.A(G299), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n841), .A2(KEYINPUT69), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n496), .A2(new_n483), .A3(new_n487), .A4(new_n498), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n954), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT56), .B(G2072), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n500), .A2(new_n984), .A3(new_n985), .A4(new_n976), .ZN(new_n986));
  INV_X1    g561(.A(new_n954), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n841), .A2(new_n976), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT112), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n841), .A2(new_n990), .A3(new_n976), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(KEYINPUT50), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n975), .A2(new_n985), .A3(new_n976), .A4(new_n977), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n986), .A2(new_n987), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT119), .B(G1956), .Z(new_n996));
  AOI211_X1 g571(.A(new_n974), .B(new_n983), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n974), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(new_n996), .ZN(new_n999));
  INV_X1    g574(.A(new_n983), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n971), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n998), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT121), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(KEYINPUT61), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT61), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n997), .B2(new_n1001), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n989), .A2(new_n991), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n987), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2067), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n954), .B1(new_n1008), .B2(new_n985), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n978), .A2(new_n1014), .A3(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1348), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1018), .A2(KEYINPUT60), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1018), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n601), .B1(new_n1018), .B2(KEYINPUT60), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n987), .B1(new_n988), .B2(new_n979), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n979), .B2(new_n978), .ZN(new_n1024));
  INV_X1    g599(.A(G1996), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT58), .B(G1341), .Z(new_n1027));
  NAND2_X1  g602(.A1(new_n1009), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n545), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n1029), .B(KEYINPUT59), .Z(new_n1030));
  NAND4_X1  g605(.A1(new_n1005), .A2(new_n1007), .A3(new_n1022), .A4(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n997), .A2(new_n1018), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1001), .B1(new_n1032), .B2(new_n591), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1031), .A2(KEYINPUT122), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT122), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT53), .B1(new_n1024), .B2(new_n802), .ZN(new_n1037));
  INV_X1    g612(.A(G1961), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(new_n1016), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT124), .B(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n953), .A2(KEYINPUT53), .A3(new_n981), .A4(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(KEYINPUT125), .A3(G301), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1016), .A2(new_n1038), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1037), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n976), .A4(new_n977), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n987), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1047), .A2(KEYINPUT53), .A3(new_n802), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1043), .B1(new_n1052), .B2(G171), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1039), .A2(G301), .A3(new_n1041), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1036), .B(new_n1042), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(G301), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1039), .A2(G171), .A3(new_n1041), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(KEYINPUT54), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1011), .A2(new_n1013), .A3(new_n1060), .A4(new_n1015), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n772), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(G168), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1063), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT51), .B1(new_n1066), .B2(KEYINPUT123), .ZN(new_n1067));
  AOI21_X1  g642(.A(G168), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1008), .B2(new_n987), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n679), .A2(G1976), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n679), .A2(G1976), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1074), .A2(KEYINPUT116), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G305), .A2(G1981), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT117), .B(G86), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n524), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n572), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(G1981), .B2(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1071), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1073), .B2(KEYINPUT52), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1073), .A2(KEYINPUT52), .A3(new_n1076), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1078), .B(new_n1086), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G303), .A2(G8), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1096), .B(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1024), .A2(G1971), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n995), .B2(G2090), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1016), .B2(G2090), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(new_n1105), .A3(G8), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1091), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1059), .A2(new_n1070), .A3(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1034), .A2(new_n1035), .A3(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1086), .A2(new_n684), .A3(new_n679), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1071), .B1(new_n1110), .B2(new_n1079), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1106), .B2(new_n1090), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1066), .A2(G168), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1091), .A2(new_n1104), .A3(new_n1106), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1100), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1091), .A2(new_n1118), .A3(new_n1106), .A4(new_n1113), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1112), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(G301), .B1(new_n1039), .B2(new_n1051), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1107), .B(new_n1121), .C1(new_n1070), .C2(KEYINPUT62), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n970), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n722), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n963), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT46), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n959), .A2(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n959), .A2(KEYINPUT126), .A3(KEYINPUT46), .A4(new_n1025), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n957), .A2(G1996), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT47), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n958), .B(KEYINPUT48), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n969), .ZN(new_n1136));
  INV_X1    g711(.A(new_n968), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n965), .A2(new_n1137), .B1(G2067), .B2(new_n740), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n959), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT127), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1125), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g717(.A(G401), .B1(new_n862), .B2(new_n869), .ZN(new_n1144));
  INV_X1    g718(.A(G227), .ZN(new_n1145));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g720(.A(G319), .B(new_n666), .C1(new_n947), .C2(new_n948), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1147), .ZN(G308));
  INV_X1    g722(.A(new_n948), .ZN(new_n1149));
  AOI21_X1  g723(.A(new_n458), .B1(new_n1149), .B2(new_n946), .ZN(new_n1150));
  NAND4_X1  g724(.A1(new_n1150), .A2(new_n1145), .A3(new_n666), .A4(new_n1144), .ZN(G225));
endmodule


