//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT81), .B1(new_n207), .B2(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(G148gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n207), .A2(G141gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n202), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G155gat), .B(G162gat), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n215), .B1(new_n214), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  INV_X1    g022(.A(G113gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G120gat), .ZN(new_n225));
  INV_X1    g024(.A(G120gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G113gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G127gat), .ZN(new_n229));
  INV_X1    g028(.A(G134gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT69), .B(G127gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n228), .B(new_n231), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g034(.A1(G127gat), .A2(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(KEYINPUT70), .A3(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n214), .A2(new_n219), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n233), .A2(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n243), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n214), .A2(KEYINPUT84), .A3(new_n219), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT84), .B1(new_n214), .B2(new_n219), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n250), .B(KEYINPUT4), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n220), .ZN(new_n258));
  INV_X1    g057(.A(new_n221), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n250), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n214), .A2(new_n219), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n242), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n249), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(KEYINPUT5), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G57gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(G85gat), .Z(new_n268));
  NOR2_X1   g067(.A1(new_n254), .A2(new_n255), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n252), .B1(new_n269), .B2(new_n242), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n247), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n264), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(new_n264), .B2(new_n273), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT6), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n277), .B(new_n268), .C1(new_n264), .C2(new_n273), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT24), .ZN(new_n296));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT66), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n300), .B(new_n294), .C1(new_n296), .C2(new_n297), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(KEYINPUT64), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n283), .A2(new_n285), .A3(new_n288), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n305), .B(new_n294), .C1(new_n296), .C2(new_n297), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n292), .A2(new_n302), .B1(new_n307), .B2(new_n290), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT27), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  AND4_X1   g112(.A1(KEYINPUT28), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n313), .B(new_n315), .C1(new_n316), .C2(KEYINPUT67), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n295), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n282), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n285), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n320), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n280), .B(new_n281), .C1(new_n308), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n290), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n286), .A2(new_n288), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n283), .A2(new_n285), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n290), .B1(new_n331), .B2(KEYINPUT65), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n330), .A2(new_n332), .A3(new_n299), .A4(new_n301), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n312), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n336));
  AOI21_X1  g135(.A(G190gat), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n318), .B1(new_n337), .B2(new_n315), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n295), .B(new_n325), .C1(new_n338), .C2(new_n314), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n334), .A2(new_n339), .A3(G226gat), .A4(G233gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n328), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343));
  INV_X1    g142(.A(G211gat), .ZN(new_n344));
  INV_X1    g143(.A(G218gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n342), .A3(new_n346), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n354), .A3(new_n340), .ZN(new_n355));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(G64gat), .ZN(new_n357));
  INV_X1    g156(.A(G92gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT80), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n353), .A2(new_n363), .A3(new_n355), .A4(new_n360), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT30), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n328), .A2(new_n354), .A3(new_n340), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n354), .B1(new_n328), .B2(new_n340), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT30), .A4(new_n360), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n355), .A4(new_n360), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n359), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n365), .B1(new_n375), .B2(KEYINPUT79), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n279), .B(new_n376), .C1(KEYINPUT79), .C2(new_n375), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n352), .A2(new_n280), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n258), .A2(new_n259), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n352), .B1(new_n246), .B2(new_n280), .ZN(new_n381));
  OAI211_X1 g180(.A(G228gat), .B(G233gat), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n245), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n269), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G228gat), .A2(G233gat), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n243), .B2(new_n245), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n384), .B(new_n385), .C1(new_n352), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n382), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(KEYINPUT86), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT85), .B(G50gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT31), .ZN(new_n394));
  XOR2_X1   g193(.A(G78gat), .B(G106gat), .Z(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n390), .B1(new_n382), .B2(new_n387), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n392), .A3(new_n397), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n334), .A2(new_n250), .A3(new_n339), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n242), .B1(new_n308), .B2(new_n327), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT71), .A4(new_n250), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G71gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G99gat), .ZN(new_n416));
  INV_X1    g215(.A(G71gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n414), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G99gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT72), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT33), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT72), .B1(new_n416), .B2(new_n420), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT32), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT73), .B1(new_n413), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n428), .B(new_n425), .C1(new_n410), .C2(new_n412), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n407), .A2(new_n408), .A3(new_n411), .A4(new_n409), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(KEYINPUT34), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(KEYINPUT34), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT32), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT33), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n413), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n421), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n430), .A2(new_n435), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n413), .A2(new_n426), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n428), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n413), .A2(KEYINPUT73), .A3(new_n426), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n435), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n404), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT35), .B1(new_n377), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n362), .A2(new_n364), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT87), .B1(new_n375), .B2(new_n365), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n398), .A2(new_n403), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n276), .A2(new_n278), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT35), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT77), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n421), .B1(new_n413), .B2(new_n437), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n464), .A2(new_n427), .A3(new_n429), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n433), .A2(new_n434), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n445), .A2(KEYINPUT77), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n466), .A2(new_n440), .A3(new_n443), .A4(new_n444), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT76), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n430), .A2(KEYINPUT76), .A3(new_n466), .A4(new_n440), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n449), .B1(new_n462), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n247), .A2(new_n270), .A3(new_n271), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n249), .ZN(new_n479));
  OR3_X1    g278(.A1(new_n260), .A2(new_n249), .A3(new_n262), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT39), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n249), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n268), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n275), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n481), .A2(KEYINPUT40), .A3(new_n268), .A4(new_n483), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT89), .B1(new_n457), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  AOI211_X1 g291(.A(new_n492), .B(new_n489), .C1(new_n455), .C2(new_n456), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n367), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n367), .A2(new_n494), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n355), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT37), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT38), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n373), .A2(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n498), .A2(new_n499), .A3(new_n359), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n460), .A2(new_n502), .A3(new_n451), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n360), .B1(new_n373), .B2(KEYINPUT37), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n404), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n491), .A2(new_n493), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n377), .A2(new_n459), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n447), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT75), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n447), .A2(new_n514), .A3(KEYINPUT36), .A4(new_n441), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT36), .B1(new_n470), .B2(new_n475), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n477), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT97), .B(G85gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n520), .A2(new_n358), .B1(KEYINPUT8), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G99gat), .B(G106gat), .Z(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(G71gat), .A2(G78gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT95), .ZN(new_n531));
  NAND2_X1  g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(KEYINPUT96), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(KEYINPUT96), .B2(KEYINPUT9), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n532), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n526), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n523), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT101), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT99), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n544), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n527), .B(KEYINPUT98), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT101), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n529), .A2(new_n552), .A3(new_n542), .A4(new_n544), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n546), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n544), .B(KEYINPUT99), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(KEYINPUT10), .A3(new_n542), .A4(new_n529), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n546), .A2(new_n550), .A3(new_n553), .ZN(new_n560));
  INV_X1    g359(.A(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G176gat), .B(G204gat), .Z(new_n563));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n559), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n559), .B2(new_n562), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n519), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(G155gat), .B(G183gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n542), .A2(KEYINPUT21), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G127gat), .ZN(new_n579));
  INV_X1    g378(.A(G8gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G15gat), .B(G22gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT16), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(G1gat), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n580), .B1(new_n583), .B2(KEYINPUT93), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(G1gat), .B2(new_n581), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(KEYINPUT21), .B2(new_n542), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n578), .B(new_n229), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n587), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n577), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n344), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n591), .A3(new_n577), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  INV_X1    g397(.A(new_n596), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G43gat), .B(G50gat), .Z(new_n602));
  NOR2_X1   g401(.A1(G29gat), .A2(G36gat), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n603), .A2(KEYINPUT14), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  INV_X1    g404(.A(G29gat), .ZN(new_n606));
  INV_X1    g405(.A(G36gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT15), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n608), .A2(new_n605), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n604), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n602), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n602), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT17), .B1(new_n619), .B2(new_n614), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n618), .B(new_n620), .C1(new_n548), .C2(new_n549), .ZN(new_n621));
  AND3_X1   g420(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(new_n614), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n555), .A2(new_n624), .A3(new_n529), .ZN(new_n625));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT100), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n621), .A2(new_n623), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n625), .A2(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n623), .A4(new_n621), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n627), .A2(KEYINPUT100), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n631), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n631), .B2(new_n634), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n601), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n586), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n620), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n586), .ZN(new_n645));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n624), .B(new_n586), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n646), .B(KEYINPUT13), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n644), .A2(KEYINPUT18), .A3(new_n645), .A4(new_n646), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G169gat), .B(G197gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G113gat), .B(G141gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT12), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT94), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n649), .A2(new_n660), .A3(new_n652), .A4(new_n653), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(KEYINPUT94), .A3(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n642), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n573), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n460), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g470(.A1(new_n573), .A2(new_n668), .A3(new_n457), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n673), .A2(new_n582), .A3(KEYINPUT42), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n582), .B1(new_n673), .B2(KEYINPUT42), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n580), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  INV_X1    g477(.A(new_n476), .ZN(new_n679));
  AOI21_X1  g478(.A(G15gat), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n516), .A2(new_n517), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n669), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n669), .A2(new_n459), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  AND2_X1   g485(.A1(new_n519), .A2(new_n640), .ZN(new_n687));
  INV_X1    g486(.A(new_n572), .ZN(new_n688));
  INV_X1    g487(.A(new_n601), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n688), .A2(new_n689), .A3(new_n667), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n691), .A2(KEYINPUT106), .A3(new_n606), .A4(new_n460), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(new_n606), .A3(new_n690), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n279), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n696));
  AND3_X1   g495(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n519), .A2(KEYINPUT107), .A3(new_n640), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n519), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n640), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n460), .A3(new_n690), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n704), .A2(KEYINPUT108), .A3(new_n460), .A4(new_n690), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(G29gat), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n691), .A2(new_n607), .A3(new_n457), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  AND3_X1   g511(.A1(new_n704), .A2(new_n457), .A3(new_n690), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n607), .B2(new_n713), .ZN(G1329gat));
  NAND4_X1  g513(.A1(new_n702), .A2(new_n681), .A3(new_n703), .A4(new_n690), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G43gat), .ZN(new_n716));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n691), .A2(new_n717), .A3(new_n679), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT47), .Z(G1330gat));
  NAND4_X1  g519(.A1(new_n704), .A2(G50gat), .A3(new_n459), .A4(new_n690), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n691), .A2(new_n459), .ZN(new_n722));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g525(.A1(new_n667), .A2(new_n519), .A3(new_n641), .A4(new_n688), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n460), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n457), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT49), .B(G64gat), .Z(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n730), .B2(new_n732), .ZN(G1333gat));
  NAND3_X1  g532(.A1(new_n727), .A2(new_n417), .A3(new_n679), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n727), .A2(new_n681), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n417), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g536(.A1(new_n727), .A2(new_n459), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(G78gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1335gat));
  INV_X1    g539(.A(new_n667), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n689), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n572), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n704), .A2(new_n460), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n519), .A2(new_n640), .A3(new_n742), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n519), .A2(KEYINPUT51), .A3(new_n640), .A4(new_n742), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n688), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n460), .A2(new_n520), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n745), .A2(new_n520), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  NAND3_X1  g552(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n749), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n746), .A2(new_n755), .A3(new_n747), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n458), .A2(G92gat), .A3(new_n572), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n702), .A2(new_n457), .A3(new_n703), .A4(new_n744), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n751), .A2(G92gat), .A3(new_n458), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(G1337gat));
  NAND3_X1  g565(.A1(new_n704), .A2(new_n681), .A3(new_n744), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(G99gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n476), .A2(new_n768), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n751), .B2(new_n770), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n702), .A2(new_n459), .A3(new_n703), .A4(new_n744), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT113), .B(G106gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n404), .A2(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n774), .B(new_n775), .C1(new_n751), .C2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n772), .A2(new_n779), .A3(new_n773), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n572), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n754), .A2(new_n756), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n779), .B1(new_n772), .B2(new_n773), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n778), .B1(new_n784), .B2(new_n775), .ZN(G1339gat));
  NAND3_X1  g584(.A1(new_n641), .A2(new_n667), .A3(new_n572), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT115), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n641), .A2(new_n788), .A3(new_n667), .A4(new_n572), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n644), .A2(new_n645), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n792), .A2(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n659), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n664), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n554), .A2(new_n561), .A3(new_n556), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n559), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n561), .B1(new_n554), .B2(new_n556), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n568), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n796), .B1(new_n802), .B2(KEYINPUT55), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n640), .A3(new_n569), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n791), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(new_n569), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n798), .B2(new_n801), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n795), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT116), .A4(new_n640), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n804), .A2(new_n665), .A3(new_n666), .A4(new_n569), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n812), .A2(new_n808), .B1(new_n572), .B2(new_n795), .ZN(new_n813));
  INV_X1    g612(.A(new_n640), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n790), .B1(new_n816), .B2(new_n601), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n817), .A2(KEYINPUT117), .A3(new_n459), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n457), .A2(new_n279), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n817), .B2(new_n459), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n818), .A2(new_n679), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n667), .ZN(new_n822));
  INV_X1    g621(.A(new_n817), .ZN(new_n823));
  INV_X1    g622(.A(new_n448), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n819), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n224), .A3(new_n741), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n821), .B2(new_n572), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n226), .A3(new_n688), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  NOR3_X1   g630(.A1(new_n821), .A2(new_n232), .A3(new_n601), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n689), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n232), .B2(new_n833), .ZN(G1342gat));
  NOR3_X1   g633(.A1(new_n825), .A2(G134gat), .A3(new_n814), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n821), .B2(new_n814), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  NOR2_X1   g637(.A1(new_n817), .A2(new_n404), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n681), .A2(new_n279), .A3(new_n457), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n798), .A2(new_n801), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT119), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n847), .B(new_n844), .C1(new_n798), .C2(new_n801), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n812), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n572), .A2(new_n795), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n814), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n811), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n790), .B1(new_n852), .B2(new_n601), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT57), .B1(new_n853), .B2(new_n404), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n841), .A2(new_n842), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G141gat), .B1(new_n855), .B2(new_n667), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n842), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n210), .A3(new_n741), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT58), .ZN(G1344gat));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n817), .B2(new_n404), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n807), .A2(new_n809), .A3(new_n640), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n689), .B1(new_n851), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n786), .B(KEYINPUT120), .Z(new_n865));
  OAI211_X1 g664(.A(new_n840), .B(new_n459), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(KEYINPUT59), .A3(new_n688), .A4(new_n842), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n855), .A2(new_n572), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(KEYINPUT59), .ZN(new_n870));
  AOI21_X1  g669(.A(G148gat), .B1(new_n858), .B2(new_n688), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n870), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n871), .ZN(G1345gat));
  NOR3_X1   g671(.A1(new_n855), .A2(new_n203), .A3(new_n601), .ZN(new_n873));
  AOI21_X1  g672(.A(G155gat), .B1(new_n858), .B2(new_n689), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  NOR3_X1   g674(.A1(new_n855), .A2(new_n204), .A3(new_n814), .ZN(new_n876));
  AOI21_X1  g675(.A(G162gat), .B1(new_n858), .B2(new_n640), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n458), .A2(new_n460), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n818), .A2(new_n679), .A3(new_n820), .A4(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n667), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n823), .A2(new_n824), .A3(new_n879), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n667), .A2(G169gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(G1348gat));
  OAI21_X1  g683(.A(G176gat), .B1(new_n880), .B2(new_n572), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n882), .A2(G176gat), .A3(new_n572), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT121), .ZN(G1349gat));
  OAI21_X1  g687(.A(G183gat), .B1(new_n880), .B2(new_n601), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n882), .A2(new_n601), .A3(new_n335), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n880), .B2(new_n814), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n882), .A2(G190gat), .A3(new_n814), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT122), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(G1351gat));
  OAI21_X1  g698(.A(new_n879), .B1(new_n516), .B2(new_n517), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT123), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n867), .A2(new_n741), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G197gat), .ZN(new_n903));
  INV_X1    g702(.A(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n839), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n667), .A2(G197gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(G1352gat));
  NOR3_X1   g706(.A1(new_n905), .A2(G204gat), .A3(new_n572), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n910), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n867), .A2(new_n688), .A3(new_n901), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G204gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(G1353gat));
  NAND4_X1  g714(.A1(new_n862), .A2(new_n866), .A3(new_n689), .A4(new_n901), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G211gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n839), .A2(new_n344), .A3(new_n689), .A4(new_n904), .ZN(new_n919));
  OR2_X1    g718(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n920));
  NAND2_X1  g719(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n916), .A2(G211gat), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT126), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n918), .A2(new_n925), .A3(new_n919), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1354gat));
  OAI21_X1  g726(.A(new_n345), .B1(new_n905), .B2(new_n814), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n867), .A2(G218gat), .A3(new_n640), .A4(new_n901), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G1355gat));
endmodule


