//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT28), .A3(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n216), .A2(new_n223), .A3(new_n217), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n219), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n214), .A2(new_n215), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n208), .A2(G183gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n204), .A2(G190gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n215), .A2(KEYINPUT24), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(KEYINPUT23), .B2(new_n220), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n229), .A2(new_n231), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G169gat), .A3(G176gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G169gat), .ZN(new_n242));
  INV_X1    g041(.A(G176gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT23), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT25), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n204), .A2(G190gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n208), .A2(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n230), .B1(new_n249), .B2(KEYINPUT24), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n236), .A2(new_n237), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n203), .B1(new_n226), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G183gat), .B(G190gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n231), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n244), .A2(new_n235), .A3(new_n217), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n237), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n214), .A2(new_n225), .A3(new_n215), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT72), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n202), .B1(new_n252), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n226), .A2(new_n251), .ZN(new_n263));
  INV_X1    g062(.A(new_n202), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n263), .A2(KEYINPUT29), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  INV_X1    g066(.A(G218gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G211gat), .A2(G218gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT71), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n276));
  NAND2_X1  g075(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n270), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G197gat), .B(G204gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n272), .A2(new_n274), .A3(new_n278), .A4(new_n279), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n266), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G8gat), .B(G36gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT75), .ZN(new_n288));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n252), .A2(new_n292), .A3(new_n261), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n293), .A2(new_n294), .A3(new_n202), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n293), .B2(new_n202), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n263), .A2(new_n202), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n286), .B(new_n291), .C1(new_n298), .C2(new_n283), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n293), .A2(new_n202), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n297), .B1(new_n302), .B2(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n293), .A2(new_n294), .A3(new_n202), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n284), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(KEYINPUT30), .A3(new_n291), .A4(new_n286), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n283), .B1(new_n303), .B2(new_n304), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT74), .B1(new_n309), .B2(new_n285), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n286), .B(new_n311), .C1(new_n298), .C2(new_n283), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n291), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT0), .ZN(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n318));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT2), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322));
  AND2_X1   g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT78), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n321), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G155gat), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT77), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(G155gat), .B2(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(G155gat), .A3(G162gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT79), .B(G155gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT80), .B(G162gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(new_n333), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n319), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n328), .A3(new_n329), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n331), .A2(new_n342), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n318), .B1(new_n350), .B2(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n330), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n320), .ZN(new_n353));
  INV_X1    g152(.A(new_n342), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n344), .A2(new_n345), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT2), .ZN(new_n357));
  INV_X1    g156(.A(new_n349), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT81), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G127gat), .ZN(new_n364));
  INV_X1    g163(.A(G127gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G134gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(G113gat), .B2(G120gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT66), .B(G113gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G120gat), .ZN(new_n372));
  INV_X1    g171(.A(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G120gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n375), .A2(new_n369), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n370), .A2(new_n372), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n350), .B2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n370), .A2(new_n372), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n367), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT4), .B1(new_n350), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n355), .A2(new_n377), .A3(new_n359), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n379), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n362), .B2(new_n378), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n350), .A2(new_n382), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n384), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(KEYINPUT82), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n383), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n377), .B1(new_n355), .B2(new_n359), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n390), .B1(new_n400), .B2(new_n394), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n388), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n317), .B(new_n392), .C1(new_n399), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n317), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n398), .B2(new_n393), .ZN(new_n405));
  INV_X1    g204(.A(new_n392), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(KEYINPUT6), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n308), .A2(new_n313), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT90), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n281), .A2(new_n292), .A3(new_n282), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n360), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n350), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n351), .B2(new_n361), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n283), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI221_X1 g221(.A(new_n416), .B1(new_n420), .B2(new_n419), .C1(new_n417), .C2(new_n283), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(G22gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n423), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n424), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n425), .A2(new_n432), .A3(new_n424), .A4(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n377), .B1(new_n226), .B2(new_n251), .ZN(new_n437));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n259), .A2(new_n260), .A3(new_n382), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT32), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(G15gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G43gat), .ZN(new_n449));
  INV_X1    g248(.A(G15gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n447), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G43gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n442), .A2(new_n444), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n453), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT32), .B(new_n441), .C1(new_n456), .C2(new_n443), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n440), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n438), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT34), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  AOI211_X1 g262(.A(new_n439), .B(new_n463), .C1(new_n437), .C2(new_n440), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n458), .A2(new_n466), .A3(KEYINPUT69), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n465), .A2(new_n455), .A3(new_n457), .ZN(new_n468));
  INV_X1    g267(.A(new_n461), .ZN(new_n469));
  INV_X1    g268(.A(new_n464), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n455), .A2(new_n457), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT69), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n413), .B1(new_n436), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n466), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n455), .A3(new_n457), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n473), .B2(new_n476), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT90), .A3(new_n435), .A4(new_n434), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n412), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT91), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT35), .ZN(new_n485));
  INV_X1    g284(.A(new_n412), .ZN(new_n486));
  INV_X1    g285(.A(new_n472), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n436), .A2(KEYINPUT35), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n479), .A2(KEYINPUT36), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n472), .A2(KEYINPUT36), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n436), .B(KEYINPUT86), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n411), .A2(new_n299), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n306), .A2(new_n498), .A3(new_n286), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n290), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT38), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n298), .A2(new_n283), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT88), .B1(new_n266), .B2(new_n284), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n504), .B(KEYINPUT37), .C1(new_n505), .C2(new_n502), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n497), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n498), .B1(new_n310), .B2(new_n312), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT38), .B1(new_n508), .B2(new_n500), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT89), .B(KEYINPUT38), .C1(new_n508), .C2(new_n500), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n379), .A2(new_n386), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n390), .ZN(new_n517));
  OR3_X1    g316(.A1(new_n400), .A2(new_n394), .A3(new_n390), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(KEYINPUT39), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n317), .B1(new_n517), .B2(KEYINPUT39), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n407), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n519), .A2(new_n520), .A3(new_n515), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n308), .B2(new_n313), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n524), .B(new_n527), .C1(new_n308), .C2(new_n313), .ZN(new_n528));
  INV_X1    g327(.A(new_n436), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n496), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n491), .A2(new_n531), .ZN(new_n532));
  NOR3_X1   g331(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n541));
  INV_X1    g340(.A(new_n538), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT94), .B(KEYINPUT15), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n542), .A2(new_n543), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n537), .A2(new_n540), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n536), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n533), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT15), .A3(new_n538), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(KEYINPUT17), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT96), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT16), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(G1gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(G1gat), .B2(new_n552), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G8gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n545), .A2(new_n549), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n551), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n556), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n562), .A4(new_n563), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT97), .B1(new_n558), .B2(new_n556), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(new_n563), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n562), .B(KEYINPUT13), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G113gat), .B(G141gat), .Z(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT12), .Z(new_n577));
  NAND4_X1  g376(.A1(new_n566), .A2(new_n567), .A3(new_n571), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n564), .A2(new_n565), .B1(new_n570), .B2(new_n569), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT98), .A3(new_n567), .A4(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n567), .ZN(new_n584));
  INV_X1    g383(.A(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT101), .ZN(new_n590));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n594), .B2(new_n595), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT103), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n601), .A2(KEYINPUT103), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(KEYINPUT103), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n609), .A2(new_n558), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n551), .A2(new_n560), .A3(new_n608), .A4(new_n605), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT104), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT104), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n559), .B2(new_n558), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(new_n551), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n610), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(new_n610), .C1(new_n612), .C2(new_n615), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n592), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n592), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G57gat), .B(G64gat), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G71gat), .B(G78gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n608), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  INV_X1    g434(.A(new_n631), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n605), .A2(new_n636), .A3(new_n608), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n626), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI211_X1 g441(.A(KEYINPUT105), .B(new_n626), .C1(new_n638), .C2(new_n639), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n625), .B1(new_n634), .B2(new_n637), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR4_X1   g447(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n640), .ZN(new_n650));
  INV_X1    g449(.A(new_n644), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT99), .B(KEYINPUT21), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G127gat), .B(G155gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n556), .B1(KEYINPUT21), .B2(new_n631), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT100), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n660), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n624), .A2(new_n654), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n532), .A2(new_n587), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT106), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n411), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  OR2_X1    g472(.A1(new_n308), .A2(new_n313), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  AND3_X1   g474(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G8gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n671), .B2(new_n674), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n676), .ZN(G1325gat));
  NAND3_X1  g479(.A1(new_n671), .A2(new_n450), .A3(new_n472), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n671), .A2(new_n494), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n450), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n671), .A2(new_n495), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  AOI21_X1  g485(.A(new_n484), .B1(new_n481), .B2(KEYINPUT35), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n489), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n513), .A2(new_n528), .A3(new_n529), .A4(new_n526), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n688), .A2(new_n485), .B1(new_n689), .B2(new_n496), .ZN(new_n690));
  INV_X1    g489(.A(new_n587), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n623), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n621), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(new_n654), .A3(new_n667), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n411), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(G29gat), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n653), .B(KEYINPUT108), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n587), .A3(new_n668), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n690), .B2(new_n694), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n694), .B1(new_n491), .B2(new_n531), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n703), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n701), .B1(new_n713), .B2(new_n698), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n411), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(G29gat), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n716), .ZN(G1328gat));
  INV_X1    g516(.A(G36gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n712), .A2(new_n674), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(KEYINPUT111), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(KEYINPUT111), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n308), .A2(new_n313), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n697), .A2(G36gat), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(G1329gat));
  OAI21_X1  g524(.A(new_n452), .B1(new_n697), .B2(new_n487), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n494), .A2(G43gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n713), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g528(.A(G50gat), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n730), .B(new_n495), .C1(new_n697), .C2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT112), .B1(new_n692), .B2(new_n696), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n730), .B1(new_n712), .B2(new_n495), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT48), .B1(new_n732), .B2(new_n733), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n730), .B1(new_n712), .B2(new_n436), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n736), .A2(KEYINPUT48), .B1(new_n737), .B2(new_n738), .ZN(G1331gat));
  INV_X1    g538(.A(new_n702), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n740), .A2(new_n691), .A3(new_n667), .A4(new_n694), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT113), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n532), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n411), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n532), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n722), .B(new_n746), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n494), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n487), .A2(G71gat), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(G71gat), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n743), .A2(new_n495), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g554(.A1(new_n691), .A2(new_n668), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT114), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n654), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n532), .A2(new_n624), .B1(new_n704), .B2(new_n705), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n694), .B(new_n709), .C1(new_n491), .C2(new_n531), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n698), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT35), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n687), .A3(new_n489), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n492), .A2(new_n493), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT86), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n436), .B(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(new_n412), .ZN(new_n769));
  INV_X1    g568(.A(new_n530), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n513), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n624), .B(new_n757), .C1(new_n765), .C2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n757), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n654), .A2(new_n594), .A3(new_n411), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n763), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NAND4_X1  g578(.A1(new_n776), .A2(new_n595), .A3(new_n674), .A4(new_n740), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n722), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n595), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT52), .ZN(G1337gat));
  OR4_X1    g582(.A1(G99gat), .A2(new_n777), .A3(new_n487), .A4(new_n653), .ZN(new_n784));
  OAI21_X1  g583(.A(G99gat), .B1(new_n762), .B2(new_n766), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n495), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n702), .A2(G106gat), .A3(new_n529), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(G106gat), .B1(new_n776), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n758), .B1(new_n707), .B2(new_n711), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n495), .ZN(new_n795));
  INV_X1    g594(.A(new_n789), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n774), .B2(new_n775), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n772), .A2(new_n773), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n708), .B2(new_n757), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n789), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n791), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n793), .B1(new_n794), .B2(new_n436), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G106gat), .B1(new_n762), .B2(new_n529), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n806), .A2(new_n807), .A3(new_n791), .A4(new_n802), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n809), .ZN(G1339gat));
  NAND2_X1  g609(.A1(new_n650), .A2(KEYINPUT105), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n638), .A2(new_n639), .A3(new_n626), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(KEYINPUT54), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n640), .A2(new_n641), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n647), .B1(new_n640), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n649), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  INV_X1    g620(.A(new_n817), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n642), .A2(new_n643), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n813), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n821), .B1(new_n824), .B2(KEYINPUT55), .ZN(new_n825));
  AND4_X1   g624(.A1(new_n821), .A2(new_n815), .A3(KEYINPUT55), .A4(new_n817), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n820), .B(new_n587), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n576), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n569), .A2(new_n570), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n583), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n654), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n624), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n624), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n668), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n691), .A2(new_n694), .A3(new_n653), .A4(new_n667), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n674), .A2(new_n698), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n495), .A2(new_n487), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n691), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n698), .B1(new_n838), .B2(new_n839), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n475), .A2(new_n480), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n722), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n691), .A2(new_n371), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT118), .ZN(G1340gat));
  NOR3_X1   g650(.A1(new_n843), .A2(new_n374), .A3(new_n702), .ZN(new_n852));
  INV_X1    g651(.A(new_n848), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n654), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n854), .B2(new_n374), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n843), .B2(new_n668), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n667), .A2(new_n365), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n848), .B2(new_n857), .ZN(G1342gat));
  NOR3_X1   g657(.A1(new_n694), .A2(G134gat), .A3(new_n674), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n847), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(KEYINPUT119), .A3(new_n861), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n843), .A2(new_n694), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT56), .B1(new_n866), .B2(G134gat), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n864), .B(new_n865), .C1(new_n867), .C2(new_n860), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n840), .A2(new_n495), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n529), .B1(new_n838), .B2(new_n839), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n766), .A2(new_n841), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT120), .Z(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G141gat), .B1(new_n876), .B2(new_n691), .ZN(new_n877));
  AND4_X1   g676(.A1(new_n722), .A2(new_n845), .A3(new_n436), .A4(new_n766), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n326), .A3(new_n587), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n882), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(G148gat), .C1(new_n876), .C2(new_n653), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n839), .B(KEYINPUT121), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n838), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n768), .A2(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n875), .A2(new_n654), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n891), .B(new_n892), .C1(new_n872), .C2(new_n871), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G148gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n887), .B1(new_n894), .B2(KEYINPUT59), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT122), .B(new_n885), .C1(new_n893), .C2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n886), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n327), .A3(new_n654), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1345gat));
  AOI21_X1  g698(.A(new_n344), .B1(new_n878), .B2(new_n667), .ZN(new_n900));
  INV_X1    g699(.A(new_n876), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n667), .A2(new_n344), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT123), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(G1346gat));
  INV_X1    g703(.A(new_n345), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n878), .A2(new_n905), .A3(new_n624), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n870), .A2(new_n624), .A3(new_n873), .A4(new_n875), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n345), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(G1347gat));
  AND4_X1   g710(.A1(new_n698), .A2(new_n840), .A3(new_n674), .A4(new_n846), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT125), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n587), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n722), .A2(new_n411), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n840), .A2(new_n842), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n691), .A2(new_n242), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n914), .A2(new_n242), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n913), .A2(new_n243), .A3(new_n654), .ZN(new_n919));
  INV_X1    g718(.A(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(G176gat), .B1(new_n920), .B2(new_n702), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1349gat));
  AOI21_X1  g721(.A(new_n204), .B1(new_n916), .B2(new_n667), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n667), .A2(new_n212), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n912), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n920), .B2(new_n694), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(KEYINPUT126), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n208), .A3(new_n624), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n930), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(G1351gat));
  NAND3_X1  g734(.A1(new_n766), .A2(new_n674), .A3(new_n436), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n411), .B(new_n936), .C1(new_n838), .C2(new_n839), .ZN(new_n937));
  INV_X1    g736(.A(G197gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n587), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT127), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n871), .A2(new_n872), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n766), .A2(new_n915), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n891), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n691), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n940), .A2(new_n945), .ZN(G1352gat));
  INV_X1    g745(.A(G204gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n937), .A2(new_n947), .A3(new_n654), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n944), .B2(new_n702), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n937), .A2(new_n267), .A3(new_n667), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n941), .A2(new_n667), .A3(new_n891), .A4(new_n943), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n944), .B2(new_n694), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n937), .A2(new_n268), .A3(new_n624), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1355gat));
endmodule


