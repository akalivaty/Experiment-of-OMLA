//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n648, new_n651, new_n652, new_n654,
    new_n655, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n462), .B2(new_n463), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(new_n463), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n462), .A2(KEYINPUT67), .A3(new_n463), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n476), .A2(G2105), .A3(new_n478), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n488), .A2(KEYINPUT69), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n474), .A2(new_n477), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n462), .B2(new_n463), .ZN(new_n498));
  AND2_X1   g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n466), .A2(G102), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n464), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n496), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(G50), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G88), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n505), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n520), .A3(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n506), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(KEYINPUT71), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n515), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n515), .A2(KEYINPUT72), .A3(new_n524), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT75), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n536), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n518), .A2(new_n520), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n543), .B1(new_n518), .B2(new_n520), .ZN(new_n545));
  OAI211_X1 g120(.A(G63), .B(G651), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n521), .A2(new_n514), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G89), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n512), .A2(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT74), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n511), .A2(new_n513), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n551), .A2(G51), .A3(G543), .A4(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n542), .A2(new_n546), .A3(new_n548), .A4(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G168));
  OAI21_X1  g131(.A(G64), .B1(new_n544), .B2(new_n545), .ZN(new_n557));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n510), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n551), .A2(G52), .A3(G543), .A4(new_n553), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n508), .A2(new_n527), .A3(G90), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n561), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n559), .B1(new_n564), .B2(new_n565), .ZN(G171));
  OAI21_X1  g141(.A(G56), .B1(new_n544), .B2(new_n545), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n510), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT77), .B(G81), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n547), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n551), .A2(G543), .A3(new_n553), .ZN(new_n572));
  INV_X1    g147(.A(G43), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  AND3_X1   g151(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G36), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G188));
  NAND4_X1  g156(.A1(new_n551), .A2(G53), .A3(G543), .A4(new_n553), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n521), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n582), .A2(new_n583), .B1(G651), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n551), .A2(G543), .A3(new_n553), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(KEYINPUT9), .A3(G53), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n547), .A2(G91), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(G299));
  NAND2_X1  g166(.A1(new_n557), .A2(new_n558), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n561), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT76), .B1(new_n560), .B2(new_n561), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(G301));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n555), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n555), .A2(new_n597), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G286));
  INV_X1    g176(.A(G166), .ZN(G303));
  NAND2_X1  g177(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n508), .A2(new_n543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(G651), .B1(new_n605), .B2(G74), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n551), .A2(G49), .A3(G543), .A4(new_n553), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n547), .A2(G87), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(G288));
  NAND3_X1  g184(.A1(new_n527), .A2(G48), .A3(G543), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n547), .A2(G86), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n510), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(G305));
  AND2_X1   g190(.A1(new_n547), .A2(G85), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n588), .A2(G47), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n605), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n618), .A2(new_n619), .A3(new_n510), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n618), .B2(new_n510), .ZN(new_n621));
  AOI211_X1 g196(.A(new_n616), .B(new_n617), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(G290));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n547), .B2(G92), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n508), .A2(new_n527), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  NOR3_X1   g202(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(G79), .A2(G543), .ZN(new_n630));
  INV_X1    g205(.A(G66), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n521), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G651), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n551), .A2(G54), .A3(G543), .A4(new_n553), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n633), .B2(new_n634), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(KEYINPUT82), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(KEYINPUT82), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n639), .A2(KEYINPUT83), .A3(new_n640), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G868), .ZN(new_n645));
  MUX2_X1   g220(.A(G301), .B(new_n644), .S(new_n645), .Z(G284));
  MUX2_X1   g221(.A(G301), .B(new_n644), .S(new_n645), .Z(G321));
  NAND2_X1  g222(.A1(G299), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n600), .B2(new_n645), .ZN(G297));
  OAI21_X1  g224(.A(new_n648), .B1(new_n600), .B2(new_n645), .ZN(G280));
  INV_X1    g225(.A(new_n644), .ZN(new_n651));
  INV_X1    g226(.A(G559), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(G860), .ZN(G148));
  OAI21_X1  g228(.A(new_n645), .B1(new_n569), .B2(new_n574), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n644), .A2(G559), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n655), .B2(new_n645), .ZN(G323));
  XNOR2_X1  g231(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g232(.A1(new_n474), .A2(new_n466), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT12), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT13), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n486), .A2(G123), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n480), .A2(G135), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n477), .A2(G111), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n465), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI221_X1 g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .C1(G99), .C2(G2105), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2096), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n669), .ZN(G156));
  XOR2_X1   g245(.A(KEYINPUT15), .B(G2435), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2438), .ZN(new_n672));
  XOR2_X1   g247(.A(G2427), .B(G2430), .Z(new_n673));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT85), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2443), .ZN(new_n678));
  XOR2_X1   g253(.A(G2451), .B(G2454), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT16), .ZN(new_n680));
  XOR2_X1   g255(.A(G1341), .B(G1348), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n678), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT86), .B(G2446), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G14), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(G401));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT88), .ZN(new_n689));
  XOR2_X1   g264(.A(G2084), .B(G2090), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(new_n691), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT17), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT18), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G2072), .A2(G2078), .ZN(new_n698));
  OAI22_X1  g273(.A1(new_n692), .A2(new_n696), .B1(new_n443), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G2096), .B(G2100), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(G227));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  XOR2_X1   g278(.A(G1961), .B(G1966), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1971), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT19), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n703), .A2(new_n704), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT89), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n709), .B1(new_n712), .B2(KEYINPUT20), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n706), .A2(new_n708), .A3(new_n710), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n713), .B(new_n714), .C1(KEYINPUT20), .C2(new_n712), .ZN(new_n715));
  XOR2_X1   g290(.A(G1991), .B(G1996), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1981), .B(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  INV_X1    g297(.A(KEYINPUT28), .ZN(new_n723));
  INV_X1    g298(.A(G26), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n486), .A2(G128), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n480), .A2(G140), .ZN(new_n728));
  NOR2_X1   g303(.A1(G104), .A2(G2105), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(new_n477), .B2(G116), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n723), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G2067), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n489), .B2(new_n490), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G35), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n736), .A2(KEYINPUT29), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(KEYINPUT29), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n738), .A2(G2090), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT101), .ZN(new_n741));
  INV_X1    g316(.A(G16), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G20), .ZN(new_n743));
  INV_X1    g318(.A(G299), .ZN(new_n744));
  OAI211_X1 g319(.A(KEYINPUT23), .B(new_n743), .C1(new_n744), .C2(new_n742), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT23), .B2(new_n743), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n740), .A2(new_n741), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G4), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n651), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1348), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n741), .B1(new_n740), .B2(new_n747), .ZN(new_n754));
  AOI21_X1  g329(.A(G2090), .B1(new_n738), .B2(new_n739), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n735), .A2(G33), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n466), .A2(G103), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  INV_X1    g333(.A(G139), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(new_n477), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n758), .B1(new_n759), .B2(new_n479), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n756), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2072), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT100), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G27), .B2(new_n735), .ZN(new_n769));
  AND3_X1   g344(.A1(new_n768), .A2(new_n735), .A3(G27), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n503), .C2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G2078), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n735), .B1(new_n774), .B2(G34), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(G34), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n472), .B2(new_n735), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n767), .B(new_n781), .C1(new_n772), .C2(new_n771), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n773), .ZN(new_n783));
  OR2_X1    g358(.A1(G29), .A2(G32), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n480), .A2(G141), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n486), .A2(G129), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n466), .A2(G105), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(new_n735), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n742), .A2(G19), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n575), .B2(new_n742), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G1341), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(G1341), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n793), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n733), .A2(G2067), .ZN(new_n800));
  NOR2_X1   g375(.A1(G5), .A2(G16), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G171), .B2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n800), .B1(G1961), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n782), .A2(new_n783), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n742), .A2(G21), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G168), .B2(new_n742), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n802), .A2(G1961), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n668), .A2(new_n735), .ZN(new_n810));
  INV_X1    g385(.A(G28), .ZN(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n811), .B2(KEYINPUT30), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(KEYINPUT30), .B2(new_n811), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT31), .B(G11), .Z(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n804), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n735), .A2(G25), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n486), .A2(G119), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n480), .A2(G131), .ZN(new_n824));
  OR2_X1    g399(.A1(G95), .A2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n822), .B1(new_n828), .B2(new_n735), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n742), .A2(G24), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n622), .B2(new_n742), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT90), .B(G1986), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n836));
  INV_X1    g411(.A(G22), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(G16), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n742), .A2(KEYINPUT93), .A3(G22), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n838), .B(new_n839), .C1(G166), .C2(new_n742), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT94), .ZN(new_n841));
  INV_X1    g416(.A(G1971), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n742), .A2(G6), .ZN(new_n844));
  INV_X1    g419(.A(G305), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(new_n742), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT32), .B(G1981), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT91), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n846), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n742), .A2(G23), .ZN(new_n851));
  INV_X1    g426(.A(G288), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n742), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT33), .B(G1976), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT92), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n853), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n843), .A2(new_n849), .A3(new_n850), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n831), .B(new_n835), .C1(new_n857), .C2(KEYINPUT34), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n860), .A2(KEYINPUT36), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n866), .A2(new_n859), .A3(new_n831), .A4(new_n835), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(KEYINPUT95), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n861), .B(KEYINPUT96), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n734), .B(new_n821), .C1(new_n864), .C2(new_n871), .ZN(G150));
  INV_X1    g447(.A(G150), .ZN(G311));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n588), .B2(G55), .ZN(new_n876));
  INV_X1    g451(.A(G67), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n603), .B2(new_n604), .ZN(new_n878));
  NAND2_X1  g453(.A1(G80), .A2(G543), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(G651), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n652), .ZN(new_n885));
  XOR2_X1   g460(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT39), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n885), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n567), .A2(new_n568), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G651), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n588), .A2(G43), .B1(new_n547), .B2(new_n570), .ZN(new_n891));
  OAI21_X1  g466(.A(G67), .B1(new_n544), .B2(new_n545), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n510), .B1(new_n892), .B2(new_n879), .ZN(new_n893));
  INV_X1    g468(.A(G55), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n572), .A2(new_n894), .B1(new_n874), .B2(new_n626), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n890), .B(new_n891), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n876), .B(new_n881), .C1(new_n569), .C2(new_n574), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n888), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n884), .B1(new_n899), .B2(G860), .ZN(G145));
  XNOR2_X1  g475(.A(new_n731), .B(new_n790), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n503), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n503), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n765), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  INV_X1    g481(.A(new_n765), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(G142), .ZN(new_n909));
  NOR2_X1   g484(.A1(G106), .A2(G2105), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(new_n477), .B2(G118), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n479), .A2(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(G130), .B2(new_n486), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n659), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n827), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n905), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n905), .B2(new_n908), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT103), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n668), .B(new_n472), .ZN(new_n919));
  XNOR2_X1  g494(.A(G162), .B(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n918), .B(new_n920), .C1(KEYINPUT103), .C2(new_n917), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n917), .B2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g501(.A1(new_n655), .A2(new_n898), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n896), .A2(new_n897), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n644), .B2(G559), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n744), .A2(new_n638), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n633), .A2(new_n634), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT81), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(G299), .A3(new_n629), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n744), .A2(new_n638), .ZN(new_n941));
  AOI21_X1  g516(.A(G299), .B1(new_n935), .B2(new_n629), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n931), .A2(new_n936), .A3(KEYINPUT41), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n927), .A2(new_n929), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n531), .A2(new_n532), .A3(G288), .ZN(new_n949));
  AOI21_X1  g524(.A(G288), .B1(new_n531), .B2(new_n532), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n845), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G166), .A2(new_n852), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n531), .A2(new_n532), .A3(G288), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(G305), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n622), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n954), .A3(new_n622), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n939), .A2(new_n959), .A3(new_n946), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n948), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n948), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(G868), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n882), .A2(new_n645), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(G295));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n964), .ZN(G331));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n555), .A2(new_n597), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n546), .A2(new_n548), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(KEYINPUT78), .A3(new_n542), .A4(new_n554), .ZN(new_n970));
  AOI21_X1  g545(.A(G301), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(G171), .A2(new_n555), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n928), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G171), .B1(new_n598), .B2(new_n599), .ZN(new_n974));
  NAND2_X1  g549(.A1(G301), .A2(G168), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n898), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n937), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n974), .A2(new_n898), .A3(new_n975), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n898), .B1(new_n974), .B2(new_n975), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n945), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n958), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n938), .B1(new_n978), .B2(new_n979), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n973), .A2(new_n943), .A3(new_n944), .A4(new_n976), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n951), .A2(new_n954), .A3(new_n622), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n955), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n985), .B2(new_n987), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n924), .B(new_n982), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n967), .B1(new_n991), .B2(KEYINPUT43), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT104), .B1(new_n981), .B2(new_n958), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(KEYINPUT105), .A3(new_n996), .A4(new_n982), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n991), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n1004));
  INV_X1    g579(.A(new_n999), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT107), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(G397));
  NAND3_X1  g587(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT108), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n467), .A2(new_n471), .A3(new_n1015), .A4(G40), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n503), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT109), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n827), .B(new_n830), .Z(new_n1024));
  AND2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(G1996), .A3(new_n790), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n731), .B(G2067), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1996), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1026), .B(new_n1028), .C1(new_n790), .C2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n622), .B(G1986), .Z(new_n1032));
  AOI211_X1 g607(.A(new_n1025), .B(new_n1031), .C1(new_n1022), .C2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT110), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n503), .A2(new_n1035), .A3(new_n1036), .A4(new_n1018), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1019), .A2(KEYINPUT50), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n773), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1018), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n807), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1038), .A2(KEYINPUT116), .A3(new_n773), .A4(new_n1039), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT114), .B(G8), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n555), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1050), .A2(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(new_n1052), .ZN(new_n1057));
  AOI211_X1 g632(.A(KEYINPUT51), .B(new_n1053), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1054), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1059), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT124), .B1(new_n1059), .B2(KEYINPUT62), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n531), .A2(G8), .A3(new_n532), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1064), .A2(KEYINPUT113), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT113), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT112), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1069), .A3(new_n1067), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1047), .A2(new_n842), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1039), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT111), .B(G2090), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1051), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1073), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1074), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1078), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1038), .A2(new_n1086), .A3(new_n1039), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1075), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1071), .A2(new_n1088), .A3(new_n1072), .ZN(new_n1089));
  OR2_X1    g664(.A1(G305), .A2(G1981), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1019), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1046), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(new_n1051), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1090), .A2(KEYINPUT49), .A3(new_n1091), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1976), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(new_n1101), .C1(new_n1100), .C2(G288), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1096), .B(new_n1051), .C1(new_n1100), .C2(G288), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT52), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1089), .A2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1083), .A2(new_n1084), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(new_n1054), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1045), .A2(KEYINPUT119), .A3(new_n772), .A4(new_n1046), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1021), .A2(new_n772), .A3(new_n1046), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1115), .A3(KEYINPUT53), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1117));
  INV_X1    g692(.A(G1961), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1116), .A2(new_n1124), .A3(new_n1119), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1126), .A2(new_n1127), .A3(G171), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1126), .B2(G171), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1063), .B1(new_n1110), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1129), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1126), .A2(new_n1127), .A3(G171), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1134), .A2(KEYINPUT123), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1062), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1088), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1050), .A2(KEYINPUT63), .A3(new_n600), .A4(new_n1051), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1106), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1089), .A2(new_n1105), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1050), .A2(new_n600), .A3(new_n1051), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1082), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1105), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(new_n1089), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1097), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1099), .A2(new_n1100), .A3(new_n852), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1090), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1146), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1096), .A2(G2067), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1117), .B2(new_n751), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G1956), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G299), .B(KEYINPUT57), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT117), .B(G2072), .Z(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT56), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1045), .A2(new_n1046), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1155), .A2(new_n641), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1158), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n641), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT58), .B(G1341), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1096), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1047), .B2(G1996), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n575), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1171), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n575), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n641), .A2(KEYINPUT60), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n639), .A2(new_n640), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1154), .A3(new_n1179), .ZN(new_n1180));
  AND4_X1   g755(.A1(new_n1168), .A2(new_n1174), .A3(new_n1175), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1166), .A2(new_n1163), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT61), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1166), .A2(new_n1184), .A3(new_n1163), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1167), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1141), .A2(new_n1142), .A3(new_n1082), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT54), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1043), .A2(new_n1044), .A3(new_n1013), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(KEYINPUT53), .A3(new_n772), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1192), .A2(KEYINPUT122), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1193), .B(new_n1123), .C1(KEYINPUT122), .C2(new_n1192), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1190), .B1(new_n1194), .B2(G171), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1128), .A2(new_n1129), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1194), .A2(G301), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1190), .B(new_n1197), .C1(G301), .C2(new_n1126), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1189), .B(new_n1059), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1152), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1033), .B1(new_n1136), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1023), .B1(new_n790), .B2(new_n1027), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1030), .B(KEYINPUT46), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT126), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT47), .ZN(new_n1206));
  NOR4_X1   g781(.A1(G290), .A2(G1986), .A3(new_n1021), .A4(new_n1017), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT48), .ZN(new_n1208));
  OR3_X1    g783(.A1(new_n1208), .A2(new_n1031), .A3(new_n1025), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n828), .A2(new_n830), .ZN(new_n1211));
  OAI22_X1  g786(.A1(new_n1031), .A2(new_n1211), .B1(G2067), .B2(new_n731), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1210), .B1(new_n1212), .B2(new_n1023), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1212), .A2(new_n1210), .A3(new_n1023), .ZN(new_n1214));
  OAI211_X1 g789(.A(new_n1206), .B(new_n1209), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OR2_X1    g792(.A1(new_n1214), .A2(new_n1213), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1218), .A2(KEYINPUT127), .A3(new_n1209), .A4(new_n1206), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1201), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g796(.A(G401), .ZN(new_n1223));
  INV_X1    g797(.A(new_n460), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n925), .A2(new_n1224), .A3(new_n721), .ZN(new_n1225));
  INV_X1    g799(.A(G227), .ZN(new_n1226));
  OR2_X1    g800(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1227));
  AND4_X1   g801(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(G308));
  NAND4_X1  g802(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(G225));
endmodule


