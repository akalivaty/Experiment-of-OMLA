//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n467), .A2(G136), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(new_n460), .B2(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  MUX2_X1   g050(.A(G100), .B(G112), .S(G2105), .Z(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n482), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT69), .B1(new_n482), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NOR2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(new_n473), .C1(new_n487), .C2(new_n486), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n494), .A3(new_n473), .A4(new_n491), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(KEYINPUT72), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT6), .B1(new_n505), .B2(new_n507), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(G543), .ZN(new_n517));
  OAI221_X1 g092(.A(new_n504), .B1(new_n514), .B2(new_n515), .C1(new_n516), .C2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n512), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(new_n526), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n533), .A2(new_n517), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n541), .A2(new_n517), .B1(new_n514), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n507), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT74), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  AND2_X1   g129(.A1(new_n513), .A2(G65), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT76), .B(G651), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n522), .A2(G91), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n520), .A2(G49), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n522), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT77), .B1(new_n572), .B2(new_n507), .ZN(new_n573));
  OAI21_X1  g148(.A(G61), .B1(new_n499), .B2(new_n500), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(new_n577), .A3(G651), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n512), .A2(G86), .A3(new_n513), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n573), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n520), .A2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n522), .A2(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n507), .C2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(new_n522), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  INV_X1    g162(.A(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n517), .A2(new_n588), .B1(new_n589), .B2(new_n507), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  MUX2_X1   g169(.A(G301), .B(new_n593), .S(new_n594), .Z(G284));
  MUX2_X1   g170(.A(G301), .B(new_n593), .S(new_n594), .Z(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n566), .B(KEYINPUT79), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  INV_X1    g175(.A(new_n593), .ZN(new_n601));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n548), .A2(new_n594), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n594), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT11), .Z(G282));
  INV_X1    g182(.A(new_n606), .ZN(G323));
  NAND2_X1  g183(.A1(new_n467), .A2(G2104), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT13), .Z(new_n612));
  INV_X1    g187(.A(G2100), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  MUX2_X1   g190(.A(G99), .B(G111), .S(G2105), .Z(new_n616));
  AOI22_X1  g191(.A1(G123), .A2(new_n474), .B1(new_n616), .B2(G2104), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  INV_X1    g193(.A(new_n467), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n614), .A2(new_n615), .A3(new_n622), .ZN(G156));
  INV_X1    g198(.A(G14), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2430), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT82), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n624), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n635), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT18), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n642), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n642), .B1(KEYINPUT17), .B2(new_n643), .ZN(new_n648));
  INV_X1    g223(.A(new_n644), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n642), .A2(new_n644), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n643), .B1(new_n651), .B2(KEYINPUT17), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n646), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n621), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  AOI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n657), .C2(new_n661), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G16), .A2(G22), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(G166), .B2(G16), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT86), .B(G1971), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(G16), .A2(G23), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT85), .Z(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(G288), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT33), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  INV_X1    g259(.A(G305), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(G16), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT32), .B(G1981), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n683), .A2(new_n688), .A3(new_n690), .ZN(new_n693));
  OR2_X1    g268(.A1(G16), .A2(G24), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G290), .B2(new_n678), .ZN(new_n695));
  INV_X1    g270(.A(G1986), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G25), .A2(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n467), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n474), .A2(G119), .ZN(new_n700));
  MUX2_X1   g275(.A(G95), .B(G107), .S(G2105), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G2104), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n698), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n695), .A2(new_n696), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n692), .A2(new_n693), .A3(new_n697), .A4(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT36), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n678), .A2(G5), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G171), .B2(new_n678), .ZN(new_n713));
  INV_X1    g288(.A(G1961), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n678), .A2(G20), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT23), .Z(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G299), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1956), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT87), .B(G1348), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n601), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G4), .B2(G16), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n715), .B(new_n719), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n678), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n678), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1966), .ZN(new_n726));
  NOR2_X1   g301(.A1(G29), .A2(G35), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G162), .B2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2090), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n726), .B(new_n731), .C1(new_n722), .C2(new_n720), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n548), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n469), .A2(KEYINPUT25), .A3(G103), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(G139), .A2(new_n467), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G127), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n460), .B2(new_n461), .ZN(new_n744));
  AND2_X1   g319(.A1(G115), .A2(G2104), .ZN(new_n745));
  OAI21_X1  g320(.A(G2105), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n737), .B1(new_n749), .B2(new_n736), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2072), .Z(new_n751));
  MUX2_X1   g326(.A(G104), .B(G116), .S(G2105), .Z(new_n752));
  AOI22_X1  g327(.A1(G128), .A2(new_n474), .B1(new_n752), .B2(G2104), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n619), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n736), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G2067), .Z(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  NAND2_X1  g336(.A1(G164), .A2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G27), .B2(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n736), .A2(G32), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n469), .A2(G105), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n765), .B(new_n767), .C1(G129), .C2(new_n474), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n467), .A2(G141), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT90), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n736), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT27), .B(G1996), .Z(new_n773));
  OAI221_X1 g348(.A(new_n760), .B1(new_n761), .B2(new_n763), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n772), .A2(new_n773), .B1(new_n763), .B2(new_n761), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT91), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT30), .B(G28), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n736), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n736), .B2(new_n620), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G34), .ZN(new_n782));
  MUX2_X1   g357(.A(new_n782), .B(G160), .S(G29), .Z(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n775), .B(new_n785), .C1(new_n784), .C2(new_n783), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n732), .A2(new_n735), .A3(new_n751), .A4(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n711), .A2(new_n723), .A3(new_n788), .ZN(G311));
  INV_X1    g364(.A(G311), .ZN(G150));
  NAND2_X1  g365(.A1(G80), .A2(G543), .ZN(new_n791));
  INV_X1    g366(.A(G67), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n501), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n507), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n520), .A2(G55), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n522), .A2(G93), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G860), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT37), .Z(new_n801));
  INV_X1    g376(.A(new_n799), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n548), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n544), .A2(new_n547), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(new_n799), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT38), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n601), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n811));
  INV_X1    g386(.A(G860), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n810), .B2(KEYINPUT39), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n801), .B1(new_n811), .B2(new_n813), .ZN(G145));
  XNOR2_X1  g389(.A(G160), .B(new_n478), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(new_n620), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n749), .A2(new_n771), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n749), .A2(new_n771), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT69), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n473), .B2(G114), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n482), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(G126), .A2(new_n474), .B1(new_n822), .B2(new_n481), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n494), .B1(new_n467), .B2(new_n491), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n755), .ZN(new_n827));
  OR3_X1    g402(.A1(new_n817), .A2(new_n818), .A3(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(G130), .A2(new_n474), .B1(new_n467), .B2(G142), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT95), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT95), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n831), .B(new_n832), .C1(G118), .C2(new_n473), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n703), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n611), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n827), .B1(new_n817), .B2(new_n818), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n828), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT96), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n836), .B1(new_n828), .B2(new_n837), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n816), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n843));
  INV_X1    g418(.A(G37), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n816), .B(new_n838), .C1(new_n840), .C2(KEYINPUT97), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n840), .A2(KEYINPUT97), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR3_X1    g422(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n843), .B1(new_n842), .B2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n601), .A2(KEYINPUT99), .A3(new_n602), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n806), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(new_n806), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n593), .A2(G299), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n587), .A2(new_n566), .A3(new_n592), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT41), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n860), .A2(new_n862), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT100), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n857), .A2(new_n858), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G290), .B(G288), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n685), .B(G303), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT42), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n866), .A2(new_n871), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n594), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n799), .A2(G868), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(G295));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n880), .B2(new_n881), .ZN(new_n884));
  INV_X1    g459(.A(new_n879), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n878), .B1(new_n866), .B2(new_n871), .ZN(new_n886));
  OAI21_X1  g461(.A(G868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(KEYINPUT101), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  OR2_X1    g466(.A1(G168), .A2(KEYINPUT102), .ZN(new_n892));
  NAND2_X1  g467(.A1(G168), .A2(KEYINPUT102), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(G301), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(G301), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n806), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n803), .A2(new_n894), .A3(new_n895), .A4(new_n805), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n870), .A2(new_n897), .A3(new_n868), .A4(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(new_n875), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n865), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n864), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n902), .A2(new_n903), .B1(new_n897), .B2(new_n898), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n863), .B(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n897), .A2(new_n898), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n865), .A2(new_n863), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n875), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n897), .A2(new_n869), .A3(new_n898), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n844), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n875), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n844), .A4(new_n913), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n891), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n921), .B(KEYINPUT43), .C1(new_n914), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n900), .A2(new_n906), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n918), .A3(new_n844), .A4(new_n913), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n917), .A2(new_n844), .A3(new_n913), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n927), .B2(KEYINPUT43), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n920), .B1(new_n929), .B2(new_n891), .ZN(G397));
  INV_X1    g505(.A(new_n720), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n493), .A2(new_n495), .ZN(new_n934));
  AOI21_X1  g509(.A(G1384), .B1(new_n934), .B2(new_n823), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT109), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(G164), .B2(G1384), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n942), .A3(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n931), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(G2067), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n601), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n948), .A2(KEYINPUT118), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(KEYINPUT118), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT116), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n562), .B2(new_n565), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n563), .B(KEYINPUT9), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n557), .A2(new_n558), .B1(new_n522), .B2(G91), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT116), .A4(new_n560), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT57), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n565), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n959), .A3(new_n955), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n826), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n945), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n941), .B1(new_n826), .B2(new_n963), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT108), .B(G1384), .C1(new_n934), .C2(new_n823), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT50), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G1956), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n971));
  AOI21_X1  g546(.A(new_n932), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT56), .B(G2072), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n961), .B(new_n962), .C1(new_n970), .C2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n949), .A2(new_n950), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n971), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n945), .B1(new_n935), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n973), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n974), .ZN(new_n982));
  INV_X1    g557(.A(G1956), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n936), .B1(new_n940), .B2(new_n942), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(new_n965), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n952), .A2(new_n959), .A3(new_n955), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n959), .B1(new_n952), .B2(new_n955), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n982), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n961), .A2(new_n962), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n991), .A2(KEYINPUT117), .A3(new_n985), .A4(new_n982), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n977), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT120), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n967), .A2(new_n968), .A3(new_n932), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT58), .B(G1341), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n997), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n946), .A2(KEYINPUT120), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n964), .A2(new_n971), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT119), .B(G1996), .ZN(new_n1003));
  AND4_X1   g578(.A1(new_n1002), .A2(new_n945), .A3(new_n973), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT121), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(new_n1004), .C1(new_n998), .C2(new_n1000), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n548), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT122), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT59), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(KEYINPUT59), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1000), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT120), .B1(new_n946), .B2(new_n999), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1005), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1007), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1001), .A2(KEYINPUT121), .A3(new_n1005), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(new_n1010), .A3(KEYINPUT59), .A4(new_n548), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  NOR4_X1   g596(.A1(new_n944), .A2(KEYINPUT60), .A3(new_n947), .A4(new_n593), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n937), .A2(new_n938), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n943), .A3(new_n945), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n720), .ZN(new_n1025));
  INV_X1    g600(.A(new_n947), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n593), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n948), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n1028), .B2(KEYINPUT60), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT61), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n990), .A2(new_n992), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT123), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n986), .A2(new_n987), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n982), .A2(new_n985), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1035), .B2(new_n988), .ZN(new_n1036));
  AND4_X1   g611(.A1(new_n1032), .A2(new_n976), .A3(new_n988), .A4(KEYINPUT61), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1029), .B(new_n1031), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n994), .B1(new_n1021), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1024), .A2(new_n714), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT125), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1961), .B1(new_n939), .B2(new_n943), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT125), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1002), .A2(new_n761), .A3(new_n945), .A4(new_n973), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n972), .A2(KEYINPUT53), .A3(new_n761), .A4(new_n973), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G171), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n967), .B2(new_n968), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n932), .B1(new_n935), .B2(new_n978), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n761), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1047), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(new_n1043), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1052), .B1(new_n1058), .B2(G301), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n939), .A2(new_n784), .A3(new_n943), .ZN(new_n1061));
  INV_X1    g636(.A(G1966), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT45), .B1(new_n940), .B2(new_n942), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n945), .B1(new_n964), .B2(new_n971), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1065), .A3(G168), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(G286), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1068), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1074), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G303), .A2(G8), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1971), .B1(new_n972), .B2(new_n973), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n940), .A2(new_n942), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n965), .B1(new_n1080), .B2(KEYINPUT50), .ZN(new_n1081));
  INV_X1    g656(.A(G2090), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1078), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1023), .A2(new_n943), .A3(new_n1082), .A4(new_n945), .ZN(new_n1086));
  INV_X1    g661(.A(G1971), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n979), .B2(new_n980), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1078), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(G8), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n946), .A2(G8), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G305), .B2(G1981), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n577), .B1(new_n576), .B2(G651), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT77), .B(new_n507), .C1(new_n574), .C2(new_n575), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n579), .A2(new_n580), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1981), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1097), .A2(new_n1099), .A3(KEYINPUT111), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n576), .A2(G651), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT49), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1092), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT49), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n568), .A2(new_n569), .A3(G1976), .A4(new_n570), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n946), .A2(G8), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT52), .ZN(new_n1114));
  INV_X1    g689(.A(G1976), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(G288), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n946), .A2(new_n1116), .A3(G8), .A4(new_n1112), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  AND4_X1   g693(.A1(new_n1085), .A2(new_n1091), .A3(new_n1111), .A4(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1060), .A2(new_n1072), .A3(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1042), .A2(new_n1044), .A3(new_n1049), .A4(G301), .ZN(new_n1121));
  OAI21_X1  g696(.A(G171), .B1(new_n1057), .B2(new_n1043), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT126), .B1(new_n1123), .B2(new_n1052), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1125), .B(KEYINPUT54), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1039), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1085), .A2(new_n1091), .A3(new_n1111), .A4(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G168), .A2(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1091), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1084), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1133), .B(KEYINPUT63), .C1(new_n1137), .C2(new_n1090), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT113), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1138), .ZN(new_n1140));
  OAI211_X1 g715(.A(G8), .B(new_n946), .C1(new_n1109), .C2(KEYINPUT49), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1109), .A2(KEYINPUT49), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1114), .B(new_n1117), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1084), .B(new_n1078), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1140), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1135), .A2(new_n1139), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G288), .A2(G1976), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1111), .A2(new_n1149), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1150));
  OAI221_X1 g725(.A(KEYINPUT112), .B1(new_n1091), .B2(new_n1143), .C1(new_n1150), .C2(new_n1092), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1143), .A2(new_n1091), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1092), .B1(new_n1154), .B2(new_n1102), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1129), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1072), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1072), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1131), .A2(new_n1122), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1135), .A2(new_n1147), .A3(new_n1139), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1167), .A2(KEYINPUT114), .A3(new_n1156), .A4(new_n1151), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1128), .A2(new_n1158), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1002), .A2(new_n932), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n755), .B(G2067), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT107), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n771), .B(G1996), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n703), .B(new_n706), .Z(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(G290), .B(G1986), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1170), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1169), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1172), .A2(new_n771), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1170), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT46), .ZN(new_n1183));
  INV_X1    g758(.A(G1996), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1170), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1186), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1182), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT47), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n704), .A2(new_n706), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1174), .A2(new_n1190), .B1(G2067), .B2(new_n755), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1170), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1186), .A2(G1986), .A3(G290), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT48), .Z(new_n1194));
  OAI21_X1  g769(.A(new_n1194), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1189), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1180), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g772(.A1(G229), .A2(G227), .A3(new_n458), .ZN(new_n1199));
  AND2_X1   g773(.A1(new_n1199), .A2(new_n640), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n1200), .B(new_n850), .C1(new_n926), .C2(new_n928), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


