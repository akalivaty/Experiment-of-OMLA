//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G50), .B2(G226), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G68), .A2(G238), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n227), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n209), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n203), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n214), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n223), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G226), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI211_X1 g0060(.A(new_n256), .B(new_n260), .C1(new_n223), .C2(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G97), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT73), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT73), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G33), .A3(G97), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n255), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n253), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G274), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n269), .A2(new_n271), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n272), .A2(new_n273), .A3(new_n255), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G238), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n267), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT74), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n280), .A3(new_n278), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G169), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n277), .A2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G179), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n279), .A2(new_n286), .A3(G169), .A4(new_n281), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n283), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n252), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(G68), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(G77), .B1(G20), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G50), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n232), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT11), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n232), .C1(G1), .C2(new_n209), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(G68), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT75), .B1(new_n303), .B2(G68), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT12), .Z(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n288), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n279), .A2(G200), .A3(new_n281), .ZN(new_n308));
  INV_X1    g0108(.A(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n284), .A2(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n303), .A2(new_n292), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n300), .B2(new_n292), .ZN(new_n314));
  XOR2_X1   g0114(.A(new_n314), .B(KEYINPUT69), .Z(new_n315));
  INV_X1    g0115(.A(new_n201), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n209), .B1(new_n316), .B2(new_n202), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  INV_X1    g0118(.A(new_n289), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n318), .A2(new_n319), .B1(new_n320), .B2(new_n294), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n297), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT9), .ZN(new_n324));
  MUX2_X1   g0124(.A(G222), .B(G223), .S(G1698), .Z(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT3), .B(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT68), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n254), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n330), .B2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n274), .A2(G226), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n270), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G190), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n324), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT10), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n323), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT15), .B(G87), .Z(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n318), .B(KEYINPUT70), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n294), .ZN(new_n349));
  INV_X1    g0149(.A(new_n303), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n349), .A2(new_n297), .B1(new_n328), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n300), .A2(G77), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n274), .A2(G244), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G232), .A2(G1698), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(G238), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n326), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n255), .C1(G107), .C2(new_n326), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n270), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n342), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n360), .A2(G179), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n353), .A2(new_n365), .A3(new_n361), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n353), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  INV_X1    g0173(.A(new_n258), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT76), .B(G33), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G223), .B2(G1698), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n356), .A2(G226), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n255), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n274), .A2(G232), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n270), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G169), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n340), .B2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n203), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT7), .B1(new_n376), .B2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G68), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n376), .A2(KEYINPUT7), .A3(G20), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n387), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n326), .B2(G20), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT77), .B(new_n393), .C1(new_n326), .C2(G20), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(G33), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n257), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n259), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n392), .B1(new_n405), .B2(G68), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n297), .B(new_n391), .C1(new_n406), .C2(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n318), .A2(new_n303), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n300), .B2(new_n318), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n384), .A2(new_n410), .A3(KEYINPUT18), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT18), .B1(new_n384), .B2(new_n410), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n391), .A2(new_n297), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n396), .A2(new_n397), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n387), .B1(new_n417), .B2(new_n290), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n414), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n380), .A2(G190), .A3(new_n270), .A4(new_n381), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n382), .A2(G200), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n407), .A2(new_n423), .A3(new_n422), .A4(new_n409), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n413), .A2(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n312), .A2(new_n345), .A3(new_n372), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT24), .ZN(new_n432));
  INV_X1    g0232(.A(G116), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n399), .A2(G33), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n209), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT22), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n209), .A2(G87), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n260), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G107), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G20), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT23), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT3), .ZN(new_n446));
  INV_X1    g0246(.A(new_n439), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(KEYINPUT22), .A3(new_n258), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n432), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n326), .A2(new_n447), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n438), .B1(new_n436), .B2(new_n209), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT24), .A3(new_n448), .A4(new_n444), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n297), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n208), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n303), .A2(new_n455), .A3(new_n232), .A4(new_n296), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G107), .ZN(new_n458));
  OR3_X1    g0258(.A1(new_n303), .A2(KEYINPUT87), .A3(G107), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT87), .B1(new_n303), .B2(G107), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT25), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n454), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n218), .A2(new_n356), .ZN(new_n464));
  INV_X1    g0264(.A(G257), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G1698), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n446), .A2(new_n258), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G294), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(new_n375), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n255), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n268), .A2(G1), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n254), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G264), .ZN(new_n478));
  INV_X1    g0278(.A(G274), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n470), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n463), .B1(G200), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n369), .B2(new_n482), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  INV_X1    g0285(.A(G244), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n446), .A2(new_n258), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n446), .A2(new_n491), .A3(new_n258), .A4(new_n487), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n218), .B2(new_n356), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n326), .B1(G33), .B2(G283), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n255), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n476), .A2(new_n465), .B1(new_n479), .B2(new_n475), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n485), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n254), .B1(new_n493), .B2(new_n496), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n499), .ZN(new_n503));
  OAI21_X1  g0303(.A(G190), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G97), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n456), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n303), .A2(G97), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n293), .A2(G77), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n441), .A2(KEYINPUT6), .A3(G97), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(new_n441), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n205), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G20), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n508), .B(new_n513), .C1(new_n417), .C2(new_n441), .ZN(new_n514));
  AOI211_X1 g0314(.A(new_n506), .B(new_n507), .C1(new_n514), .C2(new_n297), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n481), .B(KEYINPUT79), .C1(new_n465), .C2(new_n476), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT79), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n499), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n502), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n504), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n297), .ZN(new_n523));
  INV_X1    g0323(.A(new_n506), .ZN(new_n524));
  INV_X1    g0324(.A(new_n507), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n498), .A2(new_n485), .A3(new_n500), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT80), .B1(new_n502), .B2(new_n499), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n342), .A3(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n502), .A2(new_n519), .A3(G179), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n346), .A2(new_n303), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n319), .B2(new_n505), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n446), .A2(new_n209), .A3(G68), .A4(new_n258), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(new_n266), .B2(KEYINPUT19), .ZN(new_n537));
  OR2_X1    g0337(.A1(KEYINPUT81), .A2(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(KEYINPUT81), .A2(G87), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n206), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n533), .B1(new_n541), .B2(new_n297), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n457), .A2(new_n346), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n471), .A2(G274), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n254), .B(G250), .C1(G1), .C2(new_n268), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G238), .A2(G1698), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n486), .B2(G1698), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n436), .B1(new_n376), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n545), .B(new_n546), .C1(new_n549), .C2(new_n254), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n342), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n446), .A3(new_n258), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n433), .B2(new_n375), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n255), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(new_n340), .A3(new_n545), .A4(new_n546), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n544), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n456), .A2(new_n217), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n533), .B(new_n557), .C1(new_n541), .C2(new_n297), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(G200), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n554), .A2(G190), .A3(new_n545), .A4(new_n546), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n484), .A2(new_n522), .A3(new_n532), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n482), .A2(new_n342), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n470), .A2(new_n340), .A3(new_n478), .A4(new_n481), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n463), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n465), .A2(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n446), .A2(new_n258), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT84), .ZN(new_n571));
  XNOR2_X1  g0371(.A(KEYINPUT85), .B(G303), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n260), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n446), .A2(G264), .A3(G1698), .A4(new_n258), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT84), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n446), .A2(new_n575), .A3(new_n258), .A4(new_n569), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n255), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n475), .A2(G270), .A3(new_n254), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT82), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n475), .A2(new_n581), .A3(G270), .A4(new_n254), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n481), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT83), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n481), .A3(KEYINPUT83), .A4(new_n582), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n578), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(KEYINPUT21), .A3(G169), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(new_n585), .A3(G179), .A4(new_n586), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n457), .A2(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G283), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n209), .C1(G33), .C2(new_n505), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n297), .C1(new_n209), .C2(G116), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT20), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  OAI221_X1 g0397(.A(new_n591), .B1(G116), .B2(new_n303), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n587), .A2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(new_n598), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n369), .C2(new_n587), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n587), .A2(G169), .A3(new_n598), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n599), .B(new_n602), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n564), .A2(new_n568), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n431), .A2(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n556), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n507), .B1(new_n514), .B2(new_n297), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n530), .B1(new_n612), .B2(new_n524), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(new_n563), .A3(KEYINPUT26), .A4(new_n529), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT90), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n532), .B2(new_n562), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n615), .B(new_n617), .C1(new_n532), .C2(new_n562), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n611), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n599), .B1(new_n606), .B2(new_n607), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n567), .A2(KEYINPUT88), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n463), .A2(new_n565), .A3(new_n624), .A4(new_n566), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n627), .A2(new_n564), .A3(KEYINPUT89), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n484), .A2(new_n522), .A3(new_n532), .A4(new_n563), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n603), .A2(new_n605), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT86), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n599), .A3(new_n623), .A4(new_n625), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n629), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n621), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n431), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT91), .ZN(new_n639));
  INV_X1    g0439(.A(new_n344), .ZN(new_n640));
  INV_X1    g0440(.A(new_n307), .ZN(new_n641));
  INV_X1    g0441(.A(new_n367), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n311), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n413), .B1(new_n643), .B2(new_n428), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n644), .B2(new_n339), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(G369));
  INV_X1    g0446(.A(G13), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G20), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n208), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n567), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n463), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n484), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n657), .B2(new_n567), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT92), .ZN(new_n659));
  INV_X1    g0459(.A(new_n654), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n622), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT93), .Z(new_n662));
  AOI22_X1  g0462(.A1(new_n659), .A2(new_n662), .B1(new_n626), .B2(new_n660), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n601), .A2(new_n660), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n622), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n608), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0471(.A(new_n212), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n540), .A2(new_n433), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n234), .B2(new_n674), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n637), .A2(new_n660), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT97), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT89), .B1(new_n627), .B2(new_n564), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n630), .A2(new_n629), .A3(new_n635), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n654), .B1(new_n686), .B2(new_n621), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT97), .B1(new_n687), .B2(KEYINPUT29), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n634), .A2(new_n567), .A3(new_n599), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT99), .B1(new_n690), .B2(new_n564), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT99), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n630), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT98), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n618), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(new_n614), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n697), .A3(new_n556), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n683), .A2(new_n688), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n608), .A2(new_n568), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n630), .A3(new_n660), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT96), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n609), .A2(KEYINPUT96), .A3(new_n660), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n527), .A2(new_n528), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n589), .A2(new_n550), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n470), .A4(new_n478), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n520), .A2(new_n482), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT95), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n520), .A2(KEYINPUT95), .A3(new_n482), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n340), .A3(new_n550), .A4(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n587), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n654), .B1(new_n712), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n722), .B(new_n654), .C1(new_n712), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n701), .B1(new_n707), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n700), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n679), .B1(new_n728), .B2(G1), .ZN(G364));
  NAND2_X1  g0529(.A1(new_n648), .A2(G45), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n674), .A2(G1), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n668), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G330), .B2(new_n666), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n731), .B(KEYINPUT100), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n672), .A2(new_n376), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n235), .A2(new_n268), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(new_n250), .C2(new_n268), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n212), .A2(G355), .A3(new_n326), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n738), .B(new_n739), .C1(G116), .C2(new_n212), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n232), .B1(G20), .B2(new_n342), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n209), .A2(new_n369), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n340), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n209), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G322), .A2(new_n750), .B1(new_n754), .B2(G329), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n260), .ZN(new_n756));
  INV_X1    g0556(.A(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n340), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n747), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n756), .B1(G326), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n757), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n747), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G303), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n209), .B1(new_n752), .B2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G294), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n751), .A2(new_n748), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n758), .A2(new_n751), .ZN(new_n772));
  INV_X1    g0572(.A(G317), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT33), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT33), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n751), .A2(new_n762), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n771), .B(new_n776), .C1(G283), .C2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n761), .A2(new_n765), .A3(new_n768), .A4(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n772), .A2(new_n290), .B1(new_n766), .B2(new_n505), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT101), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n538), .A2(new_n539), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n763), .A2(new_n783), .B1(new_n769), .B2(new_n328), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G58), .B2(new_n750), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n260), .B1(new_n778), .B2(G107), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n754), .A2(G159), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(KEYINPUT32), .B1(G50), .B2(new_n760), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n782), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(KEYINPUT32), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n780), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n744), .ZN(new_n792));
  INV_X1    g0592(.A(new_n743), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n746), .B(new_n792), .C1(new_n666), .C2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n734), .B1(new_n735), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT102), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  INV_X1    g0597(.A(KEYINPUT107), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n660), .B1(new_n351), .B2(new_n352), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n363), .A2(new_n364), .A3(new_n366), .A4(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(new_n371), .C2(new_n799), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n680), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n803), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n637), .A2(new_n660), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(new_n725), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n731), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n735), .B1(new_n803), .B2(new_n741), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT105), .B(G143), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n750), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n769), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G159), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n816), .B2(new_n759), .C1(new_n320), .C2(new_n772), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT106), .B(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n292), .B2(new_n763), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n376), .B1(new_n821), .B2(new_n753), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n777), .A2(new_n290), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n766), .A2(new_n222), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n759), .A2(new_n826), .B1(new_n769), .B2(new_n433), .ZN(new_n827));
  INV_X1    g0627(.A(new_n772), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT103), .B(G283), .Z(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT104), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n777), .A2(new_n217), .B1(new_n753), .B2(new_n770), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n326), .B1(new_n767), .B2(G97), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n764), .A2(G107), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G294), .B2(new_n750), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n744), .B1(new_n825), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n744), .A2(new_n741), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n810), .B(new_n838), .C1(G77), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n809), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT108), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n654), .B(new_n803), .C1(new_n686), .C2(new_n621), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n367), .A2(new_n654), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n845), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n806), .A2(KEYINPUT108), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n641), .A2(new_n654), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n307), .B(new_n311), .C1(new_n309), .C2(new_n660), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n652), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n854), .A2(new_n419), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n409), .B1(new_n855), .B2(new_n415), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n411), .A2(new_n412), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n853), .B(new_n856), .C1(new_n857), .C2(new_n428), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n384), .A2(new_n410), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n410), .A2(new_n853), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n425), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n856), .B1(new_n384), .B2(new_n853), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n425), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n849), .A2(new_n852), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n860), .B1(new_n413), .B2(new_n429), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n859), .A2(new_n860), .A3(new_n425), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(new_n861), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n867), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(KEYINPUT109), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT109), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n870), .B2(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n869), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n307), .A2(new_n654), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n857), .A2(new_n652), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n871), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n683), .A2(new_n688), .A3(new_n699), .A4(new_n431), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n645), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n887), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n707), .A2(new_n724), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n891), .A2(new_n852), .A3(new_n805), .A4(new_n881), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT40), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n803), .B1(new_n707), .B2(new_n724), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n852), .A4(new_n870), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n891), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(G330), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n725), .A2(new_n431), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n898), .A2(new_n431), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n890), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n208), .B2(new_n648), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n433), .B1(new_n512), .B2(KEYINPUT35), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n233), .C1(KEYINPUT35), .C2(new_n512), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n235), .A2(G77), .A3(new_n385), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n201), .A2(new_n290), .ZN(new_n908));
  OAI211_X1 g0708(.A(G1), .B(new_n647), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n906), .A3(new_n909), .ZN(G367));
  OR2_X1    g0710(.A1(new_n558), .A2(new_n660), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n563), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(new_n556), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n735), .B1(new_n915), .B2(new_n743), .ZN(new_n916));
  INV_X1    g0716(.A(new_n346), .ZN(new_n917));
  INV_X1    g0717(.A(new_n736), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n745), .B1(new_n212), .B2(new_n917), .C1(new_n918), .C2(new_n243), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n760), .A2(new_n811), .B1(new_n828), .B2(G159), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n920), .B1(new_n320), .B2(new_n749), .C1(new_n316), .C2(new_n769), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(G77), .B2(new_n778), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n767), .A2(G68), .ZN(new_n923));
  AOI22_X1  g0723(.A1(G58), .A2(new_n764), .B1(new_n754), .B2(G137), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n922), .A2(new_n326), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n766), .A2(new_n441), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n764), .A2(KEYINPUT46), .A3(G116), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT46), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n763), .B2(new_n433), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n927), .B(new_n929), .C1(new_n468), .C2(new_n772), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT113), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n813), .A2(new_n829), .B1(new_n778), .B2(G97), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  INV_X1    g0734(.A(new_n572), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n935), .A2(new_n749), .B1(new_n759), .B2(new_n770), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n376), .B(new_n936), .C1(G317), .C2(new_n754), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n925), .B1(new_n926), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT47), .Z(new_n940));
  INV_X1    g0740(.A(new_n744), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n916), .B(new_n919), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n522), .B(new_n532), .C1(new_n515), .C2(new_n660), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n532), .B2(new_n660), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n659), .A2(new_n662), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT42), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n532), .B1(new_n943), .B2(new_n567), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n660), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n914), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n914), .B(KEYINPUT43), .Z(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT110), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT110), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n952), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n944), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n669), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n958), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n730), .A2(G1), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n967));
  OR4_X1    g0767(.A1(new_n663), .A2(new_n944), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT45), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n663), .A2(new_n969), .A3(new_n944), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n663), .B2(new_n944), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n663), .A2(new_n944), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n968), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n669), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n973), .A2(new_n971), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n977), .A2(new_n669), .A3(new_n970), .A4(new_n968), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n659), .B(new_n667), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n662), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(new_n727), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n976), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n728), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n673), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n963), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n942), .B1(new_n962), .B2(new_n985), .ZN(G387));
  INV_X1    g0786(.A(new_n735), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n376), .B1(new_n292), .B2(new_n749), .C1(new_n318), .C2(new_n772), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n763), .A2(new_n328), .B1(new_n753), .B2(new_n320), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT115), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G68), .A2(new_n813), .B1(new_n767), .B2(new_n346), .ZN(new_n991));
  INV_X1    g0791(.A(G159), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n991), .C1(new_n992), .C2(new_n759), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n988), .B(new_n993), .C1(G97), .C2(new_n778), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G322), .A2(new_n760), .B1(new_n828), .B2(G311), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n773), .B2(new_n749), .C1(new_n935), .C2(new_n769), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT48), .ZN(new_n997));
  INV_X1    g0797(.A(new_n829), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n468), .B2(new_n763), .C1(new_n766), .C2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT49), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n777), .A2(new_n433), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n376), .B(new_n1001), .C1(G326), .C2(new_n754), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n994), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n987), .B1(new_n1003), .B2(new_n941), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n676), .B(new_n268), .C1(new_n290), .C2(new_n328), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT114), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n348), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n292), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n736), .B1(new_n268), .B2(new_n240), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n675), .A2(new_n212), .A3(new_n326), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G107), .C2(new_n212), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1004), .B1(new_n745), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n659), .B2(new_n793), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT116), .Z(new_n1015));
  INV_X1    g0815(.A(new_n963), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n980), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n673), .B1(new_n1017), .B2(new_n728), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1015), .B1(new_n1016), .B2(new_n980), .C1(new_n1018), .C2(new_n981), .ZN(G393));
  AOI21_X1  g0819(.A(new_n735), .B1(new_n959), .B2(new_n743), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n376), .B1(new_n290), .B2(new_n763), .C1(new_n316), .C2(new_n772), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G77), .B2(new_n767), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1007), .A2(new_n813), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G87), .A2(new_n778), .B1(new_n754), .B2(new_n811), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n759), .A2(new_n320), .B1(new_n749), .B2(new_n992), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n326), .B1(new_n754), .B2(G322), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n441), .B2(new_n777), .C1(new_n763), .C2(new_n998), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT118), .Z(new_n1030));
  AOI22_X1  g0830(.A1(new_n572), .A2(new_n828), .B1(new_n813), .B2(G294), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n433), .C2(new_n766), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n759), .A2(new_n773), .B1(new_n749), .B2(new_n770), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT117), .Z(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1027), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n744), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n745), .B1(new_n505), .B2(new_n212), .C1(new_n918), .C2(new_n247), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1020), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n976), .A2(new_n978), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n1016), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n981), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n674), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1041), .B1(new_n982), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  NAND3_X1  g0845(.A1(new_n894), .A2(G330), .A3(new_n852), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n843), .B(new_n845), .C1(new_n687), .C2(new_n805), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT108), .B1(new_n806), .B2(new_n847), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n852), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n884), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n883), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n698), .A2(new_n660), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n847), .B1(new_n1053), .B2(new_n803), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT119), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n850), .A2(new_n851), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n850), .B2(new_n851), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n876), .B(new_n884), .C1(new_n1054), .C2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1047), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n698), .A2(new_n660), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n845), .B1(new_n1061), .B2(new_n805), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n850), .A2(new_n851), .A3(new_n1055), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n881), .B(new_n1051), .C1(new_n1062), .C2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n884), .B1(new_n849), .B2(new_n852), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1046), .C1(new_n1067), .C2(new_n883), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1060), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1069), .A2(new_n1016), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n883), .A2(new_n742), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n201), .A2(new_n778), .B1(new_n767), .B2(G159), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT54), .B(G143), .Z(new_n1073));
  NAND2_X1  g0873(.A1(new_n813), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n816), .C2(new_n772), .ZN(new_n1075));
  INV_X1    g0875(.A(G125), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n753), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n749), .A2(new_n821), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1075), .A2(new_n260), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n763), .A2(new_n320), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(G128), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1079), .B(new_n1082), .C1(new_n1083), .C2(new_n759), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT121), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n260), .B1(new_n763), .B2(new_n217), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT122), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G77), .B2(new_n767), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n760), .A2(G283), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n749), .A2(new_n433), .B1(new_n753), .B2(new_n468), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n823), .B(new_n1090), .C1(G97), .C2(new_n813), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G107), .B2(new_n828), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n744), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n839), .A2(new_n318), .ZN(new_n1095));
  AND4_X1   g0895(.A1(new_n987), .A2(new_n1071), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1070), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n852), .B1(new_n894), .B2(G330), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n849), .B1(new_n1047), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n894), .A2(G330), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1065), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1062), .A3(new_n1046), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n888), .A2(new_n645), .A3(new_n900), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1069), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1060), .A2(new_n1068), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n673), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1097), .A2(new_n1110), .ZN(G378));
  XOR2_X1   g0911(.A(new_n1104), .B(KEYINPUT123), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n323), .A2(new_n853), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n345), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n339), .A2(new_n344), .A3(new_n1114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AND4_X1   g0923(.A1(new_n895), .A2(new_n891), .A3(new_n805), .A4(new_n852), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n870), .B1(KEYINPUT40), .B2(new_n892), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n701), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n846), .A2(new_n848), .B1(new_n851), .B2(new_n850), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1127), .A2(new_n870), .B1(new_n883), .B2(new_n884), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1123), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n897), .A2(G330), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n886), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n897), .B2(G330), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n701), .B(new_n1123), .C1(new_n893), .C2(new_n896), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n887), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1113), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1113), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT124), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1113), .A2(new_n1139), .A3(KEYINPUT124), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1138), .A2(new_n1142), .A3(new_n673), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1135), .A2(new_n963), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1123), .A2(new_n741), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n917), .A2(new_n769), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G77), .A2(new_n764), .B1(new_n828), .B2(G97), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n222), .B2(new_n777), .C1(new_n441), .C2(new_n749), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(G283), .C2(new_n754), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n376), .A2(G41), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n760), .A2(G116), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1150), .A2(new_n923), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT58), .Z(new_n1154));
  OAI22_X1  g0954(.A1(new_n759), .A2(new_n1076), .B1(new_n766), .B2(new_n320), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G132), .A2(new_n828), .B1(new_n813), .B2(G137), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1083), .B2(new_n749), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(new_n764), .C2(new_n1073), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT59), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G33), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G41), .B1(new_n754), .B2(G124), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n992), .C2(new_n777), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G41), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1162), .A2(new_n1163), .B1(G50), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n744), .B1(new_n1154), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n839), .A2(new_n316), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1146), .A2(new_n732), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1145), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1144), .A2(new_n1169), .ZN(G375));
  OAI21_X1  g0970(.A(new_n987), .B1(new_n1058), .B2(new_n742), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n840), .A2(G68), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n376), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n760), .A2(G132), .B1(new_n813), .B2(G150), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n816), .B2(new_n749), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(new_n828), .C2(new_n1073), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n754), .A2(G128), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n767), .A2(G50), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G159), .A2(new_n764), .B1(new_n778), .B2(G58), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n759), .A2(new_n468), .B1(new_n769), .B2(new_n441), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G116), .B2(new_n828), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT125), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n754), .A2(G303), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n750), .A2(G283), .B1(new_n767), .B2(new_n346), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT126), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(new_n326), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G97), .A2(new_n764), .B1(new_n778), .B2(G77), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1183), .A2(new_n1184), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n941), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1171), .A2(new_n1172), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1103), .B2(new_n963), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n984), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1108), .ZN(G381));
  NAND2_X1  g0994(.A1(new_n1145), .A2(new_n1168), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1113), .A2(new_n1139), .A3(KEYINPUT124), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT124), .B1(new_n1113), .B2(new_n1139), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1109), .A2(new_n1112), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n673), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1195), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(G378), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1044), .B(new_n942), .C1(new_n962), .C2(new_n985), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1205), .A2(G396), .A3(G393), .ZN(new_n1206));
  OR4_X1    g1006(.A1(G384), .A2(new_n1204), .A3(G381), .A4(new_n1206), .ZN(G407));
  OAI211_X1 g1007(.A(G407), .B(G213), .C1(G343), .C2(new_n1204), .ZN(G409));
  NAND2_X1  g1008(.A1(G387), .A2(G390), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(G393), .B(new_n796), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1209), .A2(new_n1205), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1209), .B2(new_n1205), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT61), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1203), .B1(new_n1144), .B2(new_n1169), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n653), .A2(G213), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1199), .A2(new_n984), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1169), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1218), .B2(G378), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .A4(KEYINPUT60), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1106), .A2(new_n673), .A3(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT60), .B1(new_n1222), .B2(new_n1104), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1192), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G384), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G384), .B(new_n1192), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1215), .A2(new_n1219), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT62), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1214), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n653), .A2(KEYINPUT127), .A3(G213), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1226), .A2(new_n1227), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1195), .B1(new_n984), .B2(new_n1199), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1237), .A2(new_n1203), .B1(G213), .B2(new_n653), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1228), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT62), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1213), .B1(new_n1231), .B2(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1200), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G378), .B1(new_n1243), .B2(new_n1195), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1244), .A2(new_n1238), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT63), .B1(new_n1247), .B2(new_n1229), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1214), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT63), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1240), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1242), .A2(new_n1252), .ZN(G405));
  AND3_X1   g1053(.A1(new_n1204), .A2(new_n1244), .A3(new_n1228), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1213), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1228), .B1(new_n1204), .B2(new_n1244), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(G402));
endmodule


