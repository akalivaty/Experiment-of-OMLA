//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G68), .B2(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n203), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n203), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n221), .A2(new_n224), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n211), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT64), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n230), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n255), .B1(new_n260), .B2(new_n251), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n264));
  OAI21_X1  g0064(.A(G33), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT71), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(G33), .C1(new_n263), .C2(new_n264), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n229), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT7), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n274), .A3(new_n229), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G68), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(G58), .B(G68), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT16), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n257), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n263), .A2(new_n264), .A3(G33), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(KEYINPUT7), .B(new_n229), .C1(new_n283), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n274), .B1(new_n290), .B2(G20), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT70), .B(KEYINPUT3), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n285), .B1(new_n292), .B2(G33), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n293), .A2(KEYINPUT72), .A3(KEYINPUT7), .A4(new_n229), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G68), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT16), .B1(new_n296), .B2(new_n279), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n262), .B1(new_n282), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n215), .A2(G1698), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G223), .A2(G1698), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n300), .A2(new_n301), .B1(new_n267), .B2(new_n204), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n305));
  INV_X1    g0105(.A(G274), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n230), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n267), .B2(new_n310), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n311), .A2(G232), .A3(new_n305), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT73), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n304), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G169), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n304), .A2(G179), .A3(new_n308), .A4(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT18), .B1(new_n298), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n279), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n226), .B1(new_n272), .B2(KEYINPUT7), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n275), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n258), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n323));
  INV_X1    g0123(.A(new_n297), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n261), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n316), .A2(new_n317), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT18), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n324), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n315), .A2(G200), .ZN(new_n331));
  XOR2_X1   g0131(.A(KEYINPUT74), .B(G190), .Z(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n315), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n330), .A2(new_n331), .A3(new_n334), .A4(new_n262), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n325), .A2(KEYINPUT17), .A3(new_n331), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n329), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n278), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n341), .A2(new_n214), .B1(new_n229), .B2(G68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n229), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n216), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n257), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n345), .B(KEYINPUT11), .Z(new_n346));
  NOR2_X1   g0146(.A1(new_n260), .A2(new_n226), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n254), .A2(new_n226), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT12), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n268), .A2(new_n285), .A3(G232), .A4(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n290), .A2(KEYINPUT68), .A3(G232), .A4(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  INV_X1    g0157(.A(G1698), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n290), .A2(G226), .A3(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n355), .A2(new_n356), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n303), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n311), .A2(new_n305), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G238), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n308), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n307), .B1(new_n360), .B2(new_n303), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n363), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n352), .B1(new_n370), .B2(G190), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G232), .A2(G1698), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n358), .A2(G238), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n290), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n268), .A2(new_n285), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n210), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT67), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(KEYINPUT67), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n303), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n362), .A2(G244), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n308), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n253), .A2(G77), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n251), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n390));
  XOR2_X1   g0190(.A(KEYINPUT15), .B(G87), .Z(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n343), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n393), .B2(new_n257), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n388), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n340), .A2(new_n373), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n362), .A2(G226), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n358), .A2(G222), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G223), .A2(G1698), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n290), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n303), .C1(G77), .C2(new_n290), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n406), .A3(new_n308), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G200), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n227), .B2(G50), .ZN(new_n410));
  INV_X1    g0210(.A(G150), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n410), .B1(new_n411), .B2(new_n341), .C1(new_n250), .C2(new_n343), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n257), .B1(new_n214), .B2(new_n254), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n214), .B2(new_n260), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT9), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n408), .B1(new_n409), .B2(new_n407), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n415), .B2(new_n414), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT10), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n407), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n414), .B1(G169), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT66), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G179), .B2(new_n407), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n386), .A2(new_n372), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n396), .B1(new_n409), .B2(new_n385), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n419), .B(new_n423), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT69), .ZN(new_n427));
  INV_X1    g0227(.A(new_n368), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n367), .B1(new_n366), .B2(new_n363), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n370), .A2(G179), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n369), .A2(new_n427), .A3(new_n433), .A4(G169), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(new_n352), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n401), .A2(new_n426), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n358), .A2(G238), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n217), .B2(new_n358), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n311), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n303), .B1(new_n306), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n205), .B1(new_n445), .B2(G1), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n439), .B1(new_n451), .B2(new_n387), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n444), .A2(new_n450), .A3(KEYINPUT78), .A4(G179), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n444), .A2(new_n450), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n391), .A2(new_n253), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n226), .A2(G20), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT19), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(new_n229), .A3(G33), .A4(G97), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G97), .A2(G107), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(new_n204), .B1(new_n357), .B2(new_n229), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n456), .B1(new_n464), .B2(new_n257), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n258), .B(new_n253), .C1(G1), .C2(new_n267), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n391), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n455), .A2(new_n398), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n454), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n465), .B1(new_n204), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g0271(.A(G200), .B1(new_n444), .B2(new_n450), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n451), .A2(G190), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n269), .B1(new_n292), .B2(G33), .ZN(new_n478));
  INV_X1    g0278(.A(new_n270), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n204), .A2(G20), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(KEYINPUT79), .A3(new_n268), .A4(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n481), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(KEYINPUT22), .A3(new_n485), .ZN(new_n486));
  NOR4_X1   g0286(.A1(new_n377), .A2(KEYINPUT22), .A3(G20), .A4(new_n204), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n229), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT23), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n490), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(KEYINPUT80), .B2(KEYINPUT23), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(new_n343), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n489), .A2(KEYINPUT24), .A3(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n257), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n467), .A2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(KEYINPUT25), .C1(new_n253), .C2(G107), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n254), .A2(new_n504), .A3(new_n210), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n205), .A2(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT82), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n207), .A2(new_n358), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n303), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  AND2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n446), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n311), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n211), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(new_n311), .A3(KEYINPUT83), .A4(G264), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n522), .A2(new_n306), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G169), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n524), .A2(KEYINPUT84), .A3(new_n525), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT84), .B1(new_n524), .B2(new_n525), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n511), .A2(new_n512), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n511), .A2(new_n512), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n533), .A2(new_n534), .A3(new_n517), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n532), .B(new_n527), .C1(new_n535), .C2(new_n311), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n529), .B1(new_n387), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n477), .B1(new_n509), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n372), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT85), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n518), .A2(new_n409), .A3(new_n526), .A4(new_n527), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n542), .A3(new_n372), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT24), .B1(new_n489), .B2(new_n495), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n497), .B(new_n494), .C1(new_n486), .C2(new_n488), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n507), .B1(new_n547), .B2(new_n257), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n254), .A2(new_n206), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n467), .A2(G97), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  AND2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(new_n461), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n229), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n341), .A2(new_n216), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT75), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT75), .ZN(new_n559));
  INV_X1    g0359(.A(new_n557), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n552), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n559), .B(new_n560), .C1(new_n563), .C2(new_n229), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n295), .B2(G107), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n550), .B(new_n551), .C1(new_n566), .C2(new_n258), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n527), .B1(new_n207), .B2(new_n523), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G283), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n217), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n290), .A2(new_n358), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n571), .B1(new_n290), .B2(G250), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n570), .B(new_n573), .C1(new_n574), .C2(new_n358), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n266), .A2(G244), .A3(new_n268), .A4(new_n270), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n569), .B1(new_n577), .B2(new_n311), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n409), .ZN(new_n579));
  INV_X1    g0379(.A(new_n575), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n571), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n568), .B1(new_n582), .B2(new_n303), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n372), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n567), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n567), .B(KEYINPUT76), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n387), .B(new_n569), .C1(new_n577), .C2(new_n311), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(KEYINPUT77), .C1(new_n583), .C2(G169), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(KEYINPUT77), .B2(new_n587), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n585), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n211), .A2(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G257), .A2(G1698), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n592), .A2(new_n593), .B1(new_n594), .B2(new_n290), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n303), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n522), .A2(new_n311), .A3(G270), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n527), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n570), .B(new_n229), .C1(G33), .C2(new_n206), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(new_n257), .C1(new_n229), .C2(G116), .ZN(new_n600));
  XOR2_X1   g0400(.A(new_n600), .B(KEYINPUT20), .Z(new_n601));
  NAND2_X1  g0401(.A1(new_n467), .A2(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n254), .A2(new_n493), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n598), .A2(G169), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n598), .A2(G200), .ZN(new_n608));
  INV_X1    g0408(.A(new_n604), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n333), .C2(new_n598), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n598), .A2(KEYINPUT21), .A3(G169), .A4(new_n604), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n598), .A2(new_n387), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n604), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n607), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n538), .A2(new_n549), .A3(new_n590), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n438), .A2(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n423), .ZN(new_n617));
  INV_X1    g0417(.A(new_n329), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n388), .A2(new_n397), .A3(new_n399), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n436), .B1(new_n373), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(new_n339), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n617), .B1(new_n621), .B2(new_n419), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n607), .A2(new_n613), .A3(new_n611), .ZN(new_n623));
  INV_X1    g0423(.A(new_n536), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(G179), .B1(new_n528), .B2(G169), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n548), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n451), .A2(new_n387), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n469), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n466), .A2(new_n204), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n456), .B(new_n629), .C1(new_n464), .C2(new_n257), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n472), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n475), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n630), .B2(new_n472), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n628), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT87), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n628), .B(new_n637), .C1(new_n633), .C2(new_n634), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n626), .A2(new_n549), .A3(new_n639), .A4(new_n590), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n589), .A2(new_n567), .ZN(new_n642));
  INV_X1    g0442(.A(new_n634), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n475), .A3(new_n632), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n637), .B1(new_n644), .B2(new_n628), .ZN(new_n645));
  INV_X1    g0445(.A(new_n638), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n641), .B(new_n642), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n628), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n454), .A2(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n586), .A2(new_n649), .A3(new_n589), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n640), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n622), .B1(new_n438), .B2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G13), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G20), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n252), .ZN(new_n657));
  XNOR2_X1  g0457(.A(KEYINPUT88), .B(KEYINPUT27), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT89), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n665), .A3(G343), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n623), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n509), .A2(new_n537), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n549), .B(new_n670), .C1(new_n548), .C2(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n509), .A2(new_n537), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(KEYINPUT90), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(KEYINPUT90), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n509), .A2(new_n537), .A3(new_n667), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n614), .B1(new_n609), .B2(new_n667), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n668), .A2(new_n604), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n623), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT91), .ZN(G399));
  INV_X1    g0488(.A(new_n222), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G1), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n461), .A2(new_n204), .A3(new_n493), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n228), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n652), .A2(new_n667), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n652), .A2(KEYINPUT92), .A3(new_n667), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n639), .A2(new_n642), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n648), .B1(new_n704), .B2(KEYINPUT26), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n640), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .A3(new_n667), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n698), .A2(KEYINPUT93), .A3(new_n700), .A4(new_n699), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n703), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n518), .A2(new_n532), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n578), .A2(new_n455), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n612), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n612), .A4(new_n712), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n598), .A2(new_n455), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n387), .A3(new_n536), .A4(new_n578), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n668), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n722), .B(new_n723), .C1(new_n615), .C2(new_n668), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n710), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n695), .B1(new_n726), .B2(G1), .ZN(G364));
  OR2_X1    g0527(.A1(new_n683), .A2(G330), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n655), .A2(new_n445), .A3(G20), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n690), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n728), .A2(new_n684), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT95), .Z(new_n736));
  NOR2_X1   g0536(.A1(new_n387), .A2(G200), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n332), .A2(G20), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n377), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n387), .A2(new_n372), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n332), .A2(G20), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n229), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n737), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n743), .A2(G326), .B1(G311), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G294), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n409), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n229), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT100), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n387), .A2(G200), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT98), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n409), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n740), .B(new_n752), .C1(G303), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n741), .A2(new_n744), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n755), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G283), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n744), .A2(new_n387), .A3(new_n372), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G329), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n757), .A2(new_n763), .A3(new_n765), .A4(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n756), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n204), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n377), .B(new_n774), .C1(G107), .C2(new_n764), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT97), .B(G159), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT32), .Z(new_n780));
  OAI22_X1  g0580(.A1(new_n738), .A2(new_n225), .B1(new_n206), .B2(new_n750), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n782), .B1(new_n214), .B2(new_n742), .C1(new_n226), .C2(new_n758), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n745), .A2(new_n216), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n772), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n230), .B1(G20), .B2(new_n398), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n271), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n689), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n248), .A2(G45), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(G45), .C2(new_n228), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n290), .A2(G355), .A3(new_n222), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(G116), .C2(new_n222), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n786), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n796), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n683), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n787), .A2(new_n798), .A3(new_n800), .A4(new_n733), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n736), .A2(new_n801), .ZN(G396));
  OAI22_X1  g0602(.A1(new_n425), .A2(new_n424), .B1(new_n396), .B2(new_n667), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n400), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n619), .A2(new_n667), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(KEYINPUT103), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT103), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n698), .A2(new_n700), .A3(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  AND4_X1   g0611(.A1(new_n590), .A2(new_n626), .A3(new_n549), .A4(new_n639), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n651), .A2(new_n647), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n667), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n725), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n724), .A2(G330), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n810), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n734), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n290), .B1(new_n756), .B2(G107), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT101), .Z(new_n821));
  INV_X1    g0621(.A(new_n764), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n204), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n769), .A2(new_n824), .B1(new_n206), .B2(new_n750), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n742), .A2(new_n594), .B1(new_n826), .B2(new_n758), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n821), .A2(new_n823), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n493), .B2(new_n745), .C1(new_n748), .C2(new_n738), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n822), .A2(new_n226), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n271), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G132), .A2(new_n770), .B1(new_n756), .B2(G50), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n225), .C2(new_n750), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT102), .Z(new_n834));
  INV_X1    g0634(.A(new_n738), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(G143), .B1(G150), .B2(new_n759), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n742), .C1(new_n745), .C2(new_n778), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  OAI21_X1  g0639(.A(new_n829), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n786), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n809), .A2(new_n794), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n786), .A2(new_n794), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n216), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n733), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n819), .A2(new_n845), .ZN(G384));
  INV_X1    g0646(.A(KEYINPUT40), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n280), .A2(new_n281), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n261), .B1(new_n323), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n661), .B(new_n850), .C1(new_n329), .C2(new_n339), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n316), .A2(new_n317), .A3(new_n662), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n335), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n298), .A2(new_n661), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n325), .A2(new_n326), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT107), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n335), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n298), .A2(new_n318), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(KEYINPUT107), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n855), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n851), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n667), .A2(new_n351), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n435), .A2(KEYINPUT106), .A3(new_n352), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT106), .B1(new_n435), .B2(new_n352), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n373), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n436), .A2(new_n668), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n809), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n724), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n847), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n873), .A2(new_n724), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT108), .B1(new_n859), .B2(new_n862), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n856), .A2(new_n335), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT37), .B1(new_n857), .B2(new_n858), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT108), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n861), .A2(KEYINPUT107), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n856), .A2(new_n335), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n883), .B2(new_n857), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n877), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n298), .B(new_n661), .C1(new_n329), .C2(new_n339), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n876), .B(KEYINPUT40), .C1(new_n864), .C2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n875), .A2(new_n888), .A3(G330), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n817), .A2(new_n437), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT109), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n875), .A2(new_n888), .A3(new_n724), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n438), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n703), .A2(new_n437), .A3(new_n708), .A4(new_n709), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n622), .ZN(new_n896));
  INV_X1    g0696(.A(new_n865), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n871), .A2(new_n872), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n814), .A2(KEYINPUT105), .A3(new_n805), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT105), .B1(new_n814), .B2(new_n805), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n899), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n887), .B2(new_n864), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n869), .A2(new_n870), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n668), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n618), .A2(new_n661), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n896), .B(new_n912), .Z(new_n913));
  XNOR2_X1  g0713(.A(new_n894), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n252), .B2(new_n656), .ZN(new_n915));
  OAI21_X1  g0715(.A(G77), .B1(new_n225), .B2(new_n226), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n228), .A2(new_n916), .B1(G50), .B2(new_n226), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n655), .ZN(new_n918));
  INV_X1    g0718(.A(new_n563), .ZN(new_n919));
  OAI211_X1 g0719(.A(G20), .B(new_n309), .C1(new_n919), .C2(KEYINPUT35), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n493), .B(new_n920), .C1(KEYINPUT35), .C2(new_n919), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(new_n918), .A3(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n743), .A2(G143), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n822), .B2(new_n216), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n745), .A2(new_n214), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n926), .A2(new_n377), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n750), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G68), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n770), .A2(G137), .B1(G150), .B2(new_n835), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n759), .A2(new_n777), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n928), .A2(new_n930), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G58), .B2(new_n756), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n929), .A2(G107), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n756), .A2(G116), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT46), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n822), .A2(new_n206), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n594), .A2(new_n738), .B1(new_n742), .B2(new_n824), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT113), .B(G317), .Z(new_n941));
  AOI22_X1  g0741(.A1(new_n770), .A2(new_n941), .B1(G283), .B2(new_n746), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n937), .A2(new_n271), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G294), .B2(new_n759), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n934), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT47), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n786), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n639), .B1(new_n630), .B2(new_n667), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n648), .A2(new_n471), .A3(new_n668), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n796), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n789), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n797), .B1(new_n222), .B2(new_n392), .C1(new_n951), .C2(new_n239), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n947), .A2(new_n733), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n567), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n590), .B1(new_n954), .B2(new_n667), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n642), .A2(new_n668), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT44), .B1(new_n679), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n676), .A2(new_n677), .A3(new_n958), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n678), .A2(new_n964), .A3(new_n957), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n960), .A2(new_n962), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n685), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n960), .B(new_n961), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(new_n686), .A3(new_n959), .A4(new_n965), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n680), .B1(new_n623), .B2(new_n668), .ZN(new_n972));
  INV_X1    g0772(.A(new_n684), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n972), .A2(new_n973), .A3(new_n676), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n973), .B1(new_n972), .B2(new_n676), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n726), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n726), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n690), .B(KEYINPUT41), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n732), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n948), .A2(new_n949), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n676), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n958), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n586), .A2(new_n589), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n957), .B2(new_n670), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT111), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n668), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n982), .B(new_n985), .C1(new_n992), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n991), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n996), .B1(new_n998), .B2(new_n989), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n984), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n685), .A2(new_n958), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n997), .A2(new_n1000), .A3(new_n685), .A4(new_n958), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n953), .B1(new_n980), .B2(new_n1005), .ZN(G387));
  OR2_X1    g0806(.A1(new_n726), .A2(new_n976), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n690), .A3(new_n977), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n789), .B1(new_n236), .B2(new_n445), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n290), .A2(new_n693), .A3(new_n222), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n250), .A2(G50), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT50), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n445), .C1(new_n226), .C2(new_n216), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1011), .B1(new_n693), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n689), .A2(new_n210), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n786), .B(new_n796), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n929), .A2(new_n391), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n250), .B2(new_n758), .C1(new_n773), .C2(new_n216), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n938), .B(new_n1019), .C1(G50), .C2(new_n835), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n746), .A2(G68), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n743), .A2(G159), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n271), .B1(new_n770), .B2(G150), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n743), .A2(G322), .B1(G303), .B2(new_n746), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n824), .B2(new_n758), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n835), .B2(new_n941), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT114), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT48), .Z(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n826), .B2(new_n750), .C1(new_n748), .C2(new_n773), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT49), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n770), .A2(G326), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n764), .A2(G116), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1032), .A2(new_n271), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1024), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n734), .B(new_n1017), .C1(new_n1037), .C2(new_n786), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n680), .A2(new_n796), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1038), .A2(new_n1039), .B1(new_n976), .B2(new_n732), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1008), .A2(new_n1040), .ZN(G393));
  OAI21_X1  g0841(.A(new_n797), .B1(new_n206), .B2(new_n222), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n244), .B2(new_n789), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n750), .A2(new_n216), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n214), .B2(new_n758), .C1(new_n250), .C2(new_n745), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1046), .B(new_n823), .C1(G143), .C2(new_n770), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n756), .A2(G68), .ZN(new_n1048));
  INV_X1    g0848(.A(G159), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n411), .A2(new_n742), .B1(new_n738), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT51), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n788), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT115), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n758), .A2(new_n594), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n824), .A2(new_n738), .B1(new_n742), .B2(new_n760), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  OAI22_X1  g0856(.A1(new_n822), .A2(new_n210), .B1(new_n748), .B2(new_n745), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n377), .B1(new_n750), .B2(new_n493), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n826), .B2(new_n773), .C1(new_n739), .C2(new_n769), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1053), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n734), .B(new_n1043), .C1(new_n1061), .C2(new_n786), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n799), .B2(new_n958), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n732), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n971), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n971), .A2(new_n977), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n691), .B1(new_n971), .B2(new_n977), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  INV_X1    g0869(.A(new_n900), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n725), .A2(new_n809), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n907), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1072), .A2(new_n1073), .B1(new_n905), .B2(new_n908), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n707), .A2(new_n667), .A3(new_n811), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n805), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n900), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n887), .A2(new_n864), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n1073), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1071), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n905), .A2(new_n908), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n814), .A2(new_n805), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT105), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n814), .A2(KEYINPUT105), .A3(new_n805), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1070), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1081), .B1(new_n1086), .B2(new_n907), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1077), .A2(new_n1078), .A3(new_n1073), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n817), .A2(new_n873), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n900), .B1(new_n817), .B2(new_n811), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1092), .A2(new_n1071), .B1(new_n901), .B2(new_n902), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1070), .B1(new_n725), .B2(new_n809), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1089), .A2(new_n1094), .A3(new_n805), .A4(new_n1075), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1096), .A2(new_n622), .A3(new_n890), .A4(new_n895), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n895), .A2(new_n622), .A3(new_n890), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1080), .A2(new_n1099), .A3(new_n1090), .A4(new_n1096), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1100), .A3(new_n690), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1081), .A2(new_n794), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n756), .A2(G150), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n377), .B(new_n1104), .C1(G50), .C2(new_n764), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n743), .A2(G128), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n770), .A2(G125), .B1(G159), .B2(new_n929), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT54), .B(G143), .Z(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1109), .A2(new_n745), .B1(new_n837), .B2(new_n758), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT116), .Z(new_n1111));
  NAND4_X1  g0911(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G132), .B2(new_n835), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n774), .B(new_n830), .C1(G116), .C2(new_n835), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n377), .B1(new_n745), .B2(new_n206), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1115), .B(new_n1044), .C1(new_n743), .C2(G283), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(new_n210), .C2(new_n758), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G294), .B2(new_n770), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n786), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1102), .A2(new_n733), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n250), .B2(new_n843), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1074), .A2(new_n1079), .A3(new_n1071), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1089), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1124), .B2(new_n732), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1101), .A2(new_n1125), .ZN(G378));
  NAND2_X1  g0926(.A1(new_n419), .A2(new_n423), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT119), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n414), .A2(new_n661), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n794), .ZN(new_n1135));
  INV_X1    g0935(.A(G132), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n758), .A2(new_n1136), .B1(new_n745), .B2(new_n837), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT118), .Z(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n411), .B2(new_n750), .C1(new_n773), .C2(new_n1109), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G125), .B2(new_n743), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n738), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n764), .A2(new_n777), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G41), .B1(new_n770), .B2(G124), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1143), .A2(new_n267), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G41), .B1(new_n480), .B2(G33), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1146), .A2(new_n1147), .B1(G50), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n773), .A2(new_n216), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n822), .A2(new_n225), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n769), .A2(new_n826), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n930), .B1(new_n742), .B2(new_n493), .C1(new_n210), .C2(new_n738), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G97), .A2(new_n759), .B1(new_n746), .B2(new_n391), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT117), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n310), .A3(new_n271), .A4(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT58), .Z(new_n1158));
  OAI21_X1  g0958(.A(new_n786), .B1(new_n1149), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n843), .A2(new_n214), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1135), .A2(new_n733), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT120), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n875), .A2(new_n888), .A3(G330), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n912), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n889), .A2(new_n909), .A3(new_n911), .A4(new_n903), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1163), .B1(new_n1171), .B2(new_n1064), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1166), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1099), .A2(new_n1100), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n690), .B1(new_n1177), .B2(KEYINPUT57), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1099), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1180), .A3(KEYINPUT57), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1173), .B1(new_n1178), .B2(new_n1182), .ZN(G375));
  INV_X1    g0983(.A(KEYINPUT124), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1070), .A2(new_n794), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n843), .A2(new_n226), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n290), .B1(new_n764), .B2(G77), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT122), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n391), .B2(new_n929), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n210), .B2(new_n745), .C1(new_n594), .C2(new_n769), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n738), .A2(new_n826), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n742), .A2(new_n748), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n773), .A2(new_n206), .B1(new_n493), .B2(new_n758), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n770), .A2(G128), .B1(G150), .B2(new_n746), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n271), .B1(new_n756), .B2(G159), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n225), .C2(new_n822), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n835), .A2(G137), .B1(new_n759), .B2(new_n1108), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1136), .B2(new_n742), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT123), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(G50), .C2(new_n929), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n786), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1185), .A2(new_n733), .A3(new_n1186), .A4(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1184), .B(new_n1203), .C1(new_n1204), .C2(new_n1064), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1064), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1203), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT124), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n895), .A2(new_n622), .A3(new_n890), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1204), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n979), .B(KEYINPUT121), .Z(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1097), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1213), .ZN(G381));
  OAI211_X1 g1014(.A(new_n1068), .B(new_n953), .C1(new_n980), .C2(new_n1005), .ZN(new_n1215));
  INV_X1    g1015(.A(G396), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1008), .A2(new_n1216), .A3(new_n1040), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1215), .A2(G384), .A3(G381), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G378), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n691), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1172), .B1(new_n1222), .B2(new_n1181), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1218), .A2(new_n1219), .A3(new_n1223), .ZN(G407));
  NOR2_X1   g1024(.A1(new_n1218), .A2(new_n663), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1219), .ZN(new_n1226));
  OAI21_X1  g1026(.A(G213), .B1(new_n1225), .B2(new_n1226), .ZN(G409));
  AOI21_X1  g1027(.A(new_n1210), .B1(new_n1124), .B2(new_n1096), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1228), .B2(new_n1171), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n690), .A3(new_n1181), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1219), .B1(new_n1230), .B2(new_n1173), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1179), .A2(new_n1180), .A3(new_n1212), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(G378), .A3(new_n1172), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1210), .A2(new_n1204), .A3(KEYINPUT60), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n690), .A3(new_n1097), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT60), .B1(new_n1210), .B2(new_n1204), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1209), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n819), .A3(new_n845), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1209), .B(G384), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G213), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(G343), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1231), .A2(new_n1233), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT61), .B1(new_n1243), .B2(KEYINPUT63), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1239), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1211), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1247), .A2(new_n690), .A3(new_n1097), .A4(new_n1234), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G384), .B1(new_n1248), .B2(new_n1209), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT125), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1238), .A2(new_n1251), .A3(new_n1239), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1242), .A2(G2897), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1240), .B2(KEYINPUT125), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1258), .A3(KEYINPUT126), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1254), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(new_n1257), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1242), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1177), .A2(new_n1212), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1219), .A2(new_n1173), .A3(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1263), .B(new_n1265), .C1(new_n1223), .C2(new_n1219), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1259), .A2(new_n1262), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1266), .B2(new_n1240), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(G390), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1217), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1216), .B1(new_n1008), .B2(new_n1040), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1273), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(KEYINPUT127), .A3(new_n1217), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(new_n1277), .A3(new_n1215), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1270), .A2(new_n1215), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1276), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1244), .A2(new_n1267), .A3(new_n1269), .A4(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT62), .B1(new_n1266), .B2(new_n1240), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1266), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1242), .B1(G375), .B2(G378), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1240), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .A4(new_n1265), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1283), .A2(new_n1284), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1280), .B1(new_n1270), .B2(new_n1215), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1279), .B2(new_n1277), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1282), .A2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(G375), .A2(G378), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1226), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1286), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1226), .A2(new_n1295), .A3(new_n1240), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1281), .ZN(G402));
endmodule


