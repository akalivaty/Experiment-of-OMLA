//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  AND2_X1   g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n202), .A2(G50), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n208), .B1(new_n210), .B2(new_n211), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0020(.A(G238), .B(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT2), .B(G226), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n225), .B(new_n228), .ZN(G358));
  XOR2_X1   g0029(.A(G87), .B(G97), .Z(new_n230));
  XOR2_X1   g0030(.A(G107), .B(G116), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G50), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(G68), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n232), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(KEYINPUT81), .ZN(new_n241));
  INV_X1    g0041(.A(G169), .ZN(new_n242));
  AND2_X1   g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND2_X1  g0043(.A1(G1), .A2(G13), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n247), .A2(new_n249), .A3(G257), .A4(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G294), .ZN(new_n251));
  OR2_X1    g0051(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n252), .A2(new_n247), .A3(new_n249), .A4(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G250), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n250), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT5), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(new_n243), .B2(new_n244), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n209), .A2(KEYINPUT65), .A3(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n245), .A2(new_n256), .B1(new_n268), .B2(G264), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(KEYINPUT5), .B2(new_n261), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n274), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT76), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n258), .A2(KEYINPUT76), .A3(new_n260), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n242), .B1(new_n269), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n256), .A2(new_n245), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n268), .A2(G264), .ZN(new_n283));
  AND4_X1   g0083(.A1(G179), .A2(new_n282), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n241), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n244), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(G87), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT22), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT22), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n288), .A2(new_n292), .A3(new_n289), .A4(G87), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT23), .B1(new_n289), .B2(G107), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT23), .ZN(new_n296));
  INV_X1    g0096(.A(G107), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n289), .A2(G33), .A3(G116), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT80), .A2(KEYINPUT24), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n295), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT80), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT24), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n294), .A2(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  AOI211_X1 g0106(.A(new_n306), .B(new_n301), .C1(new_n291), .C2(new_n293), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n287), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n309), .A2(new_n289), .A3(G1), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n297), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT25), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT67), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n287), .B(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n310), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n246), .A2(G1), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n312), .B1(new_n318), .B2(G107), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n282), .A2(new_n280), .A3(new_n283), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G169), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n269), .A2(G179), .A3(new_n280), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT81), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n285), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n287), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n289), .A2(G116), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT20), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G283), .ZN(new_n330));
  INV_X1    g0130(.A(G97), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n289), .C1(G33), .C2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n328), .A2(KEYINPUT79), .A3(new_n329), .A4(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n332), .B(new_n287), .C1(new_n289), .C2(G116), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n329), .A2(KEYINPUT79), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(KEYINPUT79), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n310), .A2(new_n287), .ZN(new_n338));
  INV_X1    g0138(.A(G116), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n317), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n309), .A2(G1), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n338), .A2(new_n340), .B1(new_n327), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n333), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n247), .A2(new_n249), .A3(G257), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n252), .A2(new_n253), .ZN(new_n346));
  INV_X1    g0146(.A(G303), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n345), .A2(new_n346), .B1(new_n288), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n245), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n263), .A2(new_n265), .A3(G270), .A4(new_n267), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n280), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n344), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(G169), .A3(new_n343), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT21), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT21), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n352), .A2(new_n357), .A3(G169), .A4(new_n343), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n325), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n287), .B(KEYINPUT67), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n310), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n274), .A2(G20), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G50), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n289), .B1(new_n201), .B2(new_n233), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT8), .B(G58), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n289), .A2(G33), .ZN(new_n367));
  INV_X1    g0167(.A(G150), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G20), .A2(G33), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n361), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n310), .A2(new_n233), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n364), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT66), .B(G1698), .Z(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G222), .A3(new_n288), .ZN(new_n377));
  INV_X1    g0177(.A(G77), .ZN(new_n378));
  INV_X1    g0178(.A(G223), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n288), .A2(G1698), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n377), .B1(new_n378), .B2(new_n288), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n245), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n243), .A2(new_n264), .A3(new_n244), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT65), .B1(new_n209), .B2(new_n266), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n383), .A2(new_n384), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n274), .B(G274), .C1(G41), .C2(G45), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n387), .A2(G226), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(G179), .ZN(new_n393));
  AOI211_X1 g0193(.A(new_n375), .B(new_n393), .C1(new_n242), .C2(new_n392), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT9), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n374), .B1(new_n392), .B2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n375), .A2(KEYINPUT9), .ZN(new_n397));
  INV_X1    g0197(.A(new_n392), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G190), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n396), .A2(new_n397), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n394), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n247), .A2(new_n249), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G107), .ZN(new_n406));
  INV_X1    g0206(.A(G238), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n406), .B1(new_n254), .B2(new_n222), .C1(new_n407), .C2(new_n380), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n245), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n387), .A2(G244), .B1(new_n388), .B2(new_n390), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G190), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT68), .ZN(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT15), .B(G87), .Z(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n367), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n366), .A2(new_n370), .B1(new_n289), .B2(new_n378), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n287), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n378), .B1(new_n274), .B2(G20), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n338), .A2(new_n420), .B1(new_n378), .B2(new_n310), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n411), .A2(G200), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n413), .B1(KEYINPUT68), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n411), .A2(G179), .ZN(new_n427));
  AOI21_X1  g0227(.A(G169), .B1(new_n409), .B2(new_n410), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n427), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n404), .A2(KEYINPUT69), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT69), .B1(new_n404), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n310), .A2(new_n235), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT12), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n369), .A2(G50), .B1(G20), .B2(new_n235), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n378), .B2(new_n367), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n361), .A2(KEYINPUT11), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n338), .A2(G68), .A3(new_n363), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n361), .A2(new_n437), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(KEYINPUT11), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G97), .ZN(new_n444));
  INV_X1    g0244(.A(G226), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n254), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n245), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n265), .A2(new_n267), .A3(G238), .A4(new_n385), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n390), .A2(new_n265), .A3(new_n267), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n412), .B1(new_n451), .B2(KEYINPUT13), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT13), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(new_n453), .A3(new_n450), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n442), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT70), .A3(new_n454), .ZN(new_n457));
  OR3_X1    g0257(.A1(new_n451), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(G200), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n458), .A3(G169), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT14), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n457), .A2(new_n458), .A3(new_n464), .A4(G169), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(G179), .A3(new_n454), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n461), .B1(new_n467), .B2(new_n442), .ZN(new_n468));
  INV_X1    g0268(.A(new_n366), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n363), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n316), .A2(new_n470), .B1(new_n315), .B2(new_n469), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT7), .B1(new_n405), .B2(new_n289), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT7), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n473), .B(G20), .C1(new_n247), .C2(new_n249), .ZN(new_n474));
  OAI21_X1  g0274(.A(G68), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G58), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n235), .ZN(new_n477));
  OAI21_X1  g0277(.A(G20), .B1(new_n477), .B2(new_n201), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n369), .A2(G159), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT16), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n326), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n475), .A2(KEYINPUT16), .A3(new_n481), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n471), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n247), .A2(new_n249), .A3(G226), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G87), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n254), .C2(new_n379), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n245), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n389), .B1(new_n386), .B2(new_n222), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n388), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n353), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n489), .A2(new_n245), .B1(new_n388), .B2(new_n491), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n242), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT18), .B1(new_n486), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n473), .B1(new_n288), .B2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n405), .A2(KEYINPUT7), .A3(new_n289), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n235), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n483), .B1(new_n501), .B2(new_n480), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n485), .A2(new_n502), .A3(new_n287), .ZN(new_n503));
  INV_X1    g0303(.A(new_n471), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n493), .A2(G169), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n495), .A2(G179), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT18), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n498), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(G190), .B1(new_n388), .B2(new_n491), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n490), .A2(KEYINPUT71), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT71), .B1(new_n490), .B2(new_n511), .ZN(new_n513));
  AOI21_X1  g0313(.A(G200), .B1(new_n490), .B2(new_n492), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n503), .A2(new_n504), .ZN(new_n516));
  NAND2_X1  g0316(.A1(KEYINPUT72), .A2(KEYINPUT17), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT72), .A2(KEYINPUT17), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n490), .A2(new_n511), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G200), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n493), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n490), .A2(KEYINPUT71), .A3(new_n511), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n521), .B1(new_n486), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT73), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n521), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n515), .B2(new_n516), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n486), .A2(new_n528), .A3(new_n517), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT73), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n510), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n433), .A2(new_n468), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  INV_X1    g0338(.A(G244), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n254), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n376), .A2(new_n288), .A3(KEYINPUT4), .A4(G244), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n247), .A2(new_n249), .A3(G250), .A4(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n330), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n245), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(new_n267), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n275), .A2(new_n276), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT76), .B1(new_n258), .B2(new_n260), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n545), .B1(new_n548), .B2(new_n272), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n544), .A2(new_n412), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n245), .B2(new_n543), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(G200), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n317), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n362), .A2(G97), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n331), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n556), .A2(new_n557), .B1(new_n297), .B2(new_n558), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n559), .A2(new_n289), .B1(new_n378), .B2(new_n370), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n297), .B1(new_n499), .B2(new_n500), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n287), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n310), .A2(new_n331), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n555), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n555), .A2(new_n562), .A3(KEYINPUT75), .A4(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n553), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n544), .A2(new_n550), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n353), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n552), .A2(new_n242), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n269), .A2(G190), .A3(new_n280), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n321), .A2(G200), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n308), .A2(new_n319), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n569), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n245), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n247), .A2(new_n249), .A3(G244), .A4(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G116), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n376), .A2(new_n288), .A3(G238), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(G250), .B1(new_n274), .B2(G45), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n270), .B2(new_n258), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n388), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n583), .A2(new_n587), .A3(new_n412), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n580), .B(new_n579), .C1(new_n254), .C2(new_n407), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n245), .B1(new_n388), .B2(new_n585), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n525), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT77), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND3_X1  g0396(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n289), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n367), .B2(new_n331), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n288), .A2(new_n289), .A3(G68), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT78), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(new_n599), .C1(new_n367), .C2(new_n331), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n287), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n416), .A2(new_n310), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n314), .A2(G87), .A3(new_n315), .A4(new_n554), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n592), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n318), .A2(new_n415), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n606), .A3(new_n607), .ZN(new_n613));
  OAI21_X1  g0413(.A(G169), .B1(new_n583), .B2(new_n587), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n590), .A2(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n343), .B1(new_n352), .B2(G200), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n412), .B2(new_n352), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n360), .A2(new_n537), .A3(new_n577), .A4(new_n622), .ZN(G372));
  AOI221_X4 g0423(.A(new_n353), .B1(new_n388), .B2(new_n585), .C1(new_n589), .C2(new_n245), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n589), .A2(new_n245), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n242), .B1(new_n625), .B2(new_n586), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT82), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT82), .B1(new_n614), .B2(new_n615), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n613), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n570), .A2(G169), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n552), .A2(G179), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n567), .A2(new_n568), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n611), .A3(new_n630), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n633), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n565), .ZN(new_n639));
  XOR2_X1   g0439(.A(KEYINPUT84), .B(KEYINPUT26), .Z(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n639), .A2(new_n617), .A3(new_n611), .A4(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n322), .A2(new_n323), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n320), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT83), .B1(new_n359), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n645), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n609), .A2(new_n588), .A3(new_n591), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n627), .B1(new_n624), .B2(new_n626), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT82), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n652), .B2(new_n613), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n647), .A2(new_n577), .A3(new_n648), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n537), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT85), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n505), .A2(new_n506), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n516), .A2(new_n508), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n508), .B1(new_n516), .B2(new_n658), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n498), .A2(new_n509), .A3(KEYINPUT85), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n467), .A2(new_n442), .B1(new_n460), .B2(new_n429), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n401), .A2(new_n403), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n394), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n656), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT86), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n341), .A2(new_n289), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n344), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n359), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n621), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n320), .A2(new_n678), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n325), .A2(new_n576), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n325), .B2(new_n679), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n359), .A2(new_n678), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n689), .A2(new_n685), .B1(new_n645), .B2(new_n678), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n688), .A2(new_n690), .ZN(G399));
  NAND3_X1  g0491(.A1(new_n595), .A2(new_n339), .A3(new_n596), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT87), .Z(new_n693));
  INV_X1    g0493(.A(new_n206), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n693), .A2(new_n274), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n211), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  OAI21_X1  g0499(.A(new_n640), .B1(new_n618), .B2(new_n573), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n635), .B2(new_n636), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n325), .A2(new_n359), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n577), .A2(new_n702), .A3(new_n653), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n703), .A3(new_n630), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .A3(new_n679), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n678), .B1(new_n643), .B2(new_n654), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT88), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n705), .B1(new_n708), .B2(KEYINPUT29), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n577), .A2(new_n360), .A3(new_n622), .A4(new_n679), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n542), .A2(new_n330), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n376), .A2(new_n288), .A3(G244), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n538), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n578), .B1(new_n715), .B2(new_n541), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n321), .B1(new_n716), .B2(new_n549), .ZN(new_n717));
  INV_X1    g0517(.A(new_n590), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n352), .A3(new_n353), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n347), .B1(new_n247), .B2(new_n249), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n247), .A2(new_n249), .A3(G257), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n376), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n578), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n351), .B1(new_n548), .B2(new_n272), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n552), .A2(new_n624), .A3(new_n727), .A4(new_n269), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n282), .A2(new_n283), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n352), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n552), .A4(new_n624), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n720), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n712), .B1(new_n734), .B2(new_n679), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n678), .A2(KEYINPUT31), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(G330), .B1(new_n711), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n709), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n699), .B1(new_n739), .B2(G1), .ZN(G364));
  INV_X1    g0540(.A(new_n695), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n309), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n274), .B1(new_n742), .B2(G45), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(KEYINPUT89), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT89), .ZN(new_n745));
  INV_X1    g0545(.A(new_n743), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n695), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n288), .A2(G355), .A3(new_n206), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n239), .A2(new_n257), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n694), .A2(new_n288), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G45), .B2(new_n211), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(G116), .B2(new_n206), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n244), .B1(G20), .B2(new_n242), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n748), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n289), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n412), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n297), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n405), .B(new_n763), .C1(G87), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT90), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n289), .A2(new_n353), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(KEYINPUT32), .B1(new_n774), .B2(G58), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(new_n525), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n412), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n289), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n775), .B1(new_n233), .B2(new_n777), .C1(new_n331), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n772), .A2(new_n412), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n772), .A2(new_n768), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n782), .A2(G68), .B1(new_n784), .B2(G77), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(KEYINPUT32), .B2(new_n771), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n774), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n788), .A2(new_n789), .B1(new_n762), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n779), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(G294), .B2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n776), .A2(G326), .B1(new_n765), .B2(G303), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n782), .A2(new_n795), .B1(new_n784), .B2(G311), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n288), .B1(new_n770), .B2(G329), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n767), .A2(new_n787), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n756), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n759), .B1(new_n760), .B2(new_n799), .C1(new_n682), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n683), .A2(new_n748), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n682), .A2(G330), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(G396));
  INV_X1    g0604(.A(new_n708), .ZN(new_n805));
  INV_X1    g0605(.A(new_n429), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n678), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n423), .A2(new_n425), .B1(new_n422), .B2(new_n679), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n806), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n805), .A2(new_n810), .B1(new_n706), .B2(new_n809), .ZN(new_n811));
  INV_X1    g0611(.A(new_n738), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(KEYINPUT94), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(KEYINPUT94), .ZN(new_n815));
  INV_X1    g0615(.A(new_n748), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n811), .B2(new_n812), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n757), .A2(new_n754), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n748), .B1(new_n378), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n782), .A2(G150), .B1(new_n784), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n821), .B1(new_n788), .B2(new_n822), .C1(new_n823), .C2(new_n777), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n288), .B1(new_n769), .B2(new_n827), .C1(new_n233), .C2(new_n764), .ZN(new_n828));
  INV_X1    g0628(.A(new_n762), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G68), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n476), .B2(new_n779), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n826), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n824), .A2(new_n825), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n782), .A2(G283), .B1(new_n784), .B2(G116), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n347), .B2(new_n777), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT91), .ZN(new_n836));
  INV_X1    g0636(.A(G87), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n762), .B1(new_n764), .B2(new_n297), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n405), .B1(new_n769), .B2(new_n839), .C1(new_n779), .C2(new_n331), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n838), .B(new_n840), .C1(G294), .C2(new_n774), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n832), .A2(new_n833), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n820), .B1(new_n760), .B2(new_n842), .C1(new_n809), .C2(new_n755), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n818), .A2(new_n843), .ZN(G384));
  NOR2_X1   g0644(.A1(new_n210), .A2(new_n339), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n559), .B(KEYINPUT95), .Z(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT35), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT36), .ZN(new_n851));
  OR3_X1    g0651(.A1(new_n211), .A2(new_n378), .A3(new_n477), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n234), .B(KEYINPUT96), .Z(new_n853));
  AOI211_X1 g0653(.A(new_n274), .B(G13), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n537), .B(new_n705), .C1(new_n708), .C2(KEYINPUT29), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n670), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n528), .A2(new_n504), .A3(new_n503), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n485), .A2(new_n502), .A3(new_n361), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n504), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n658), .ZN(new_n862));
  INV_X1    g0662(.A(new_n676), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n859), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n507), .A2(KEYINPUT97), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n516), .A2(new_n863), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n866), .B1(new_n507), .B2(KEYINPUT97), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n865), .A2(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT38), .B(new_n871), .C1(new_n536), .C2(new_n864), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n532), .A2(new_n533), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n659), .A2(new_n660), .A3(new_n657), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT85), .B1(new_n498), .B2(new_n509), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n868), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n516), .A2(new_n658), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n859), .A2(new_n880), .A3(new_n868), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT98), .ZN(new_n883));
  INV_X1    g0683(.A(new_n870), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n884), .A2(new_n859), .A3(new_n867), .A4(new_n868), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT98), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n886), .A3(KEYINPUT37), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n879), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n858), .B1(new_n873), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n871), .B1(new_n536), .B2(new_n864), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n467), .A2(new_n442), .A3(new_n679), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n663), .A2(new_n863), .ZN(new_n900));
  INV_X1    g0700(.A(new_n510), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n665), .B2(new_n666), .ZN(new_n902));
  INV_X1    g0702(.A(new_n864), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n904), .B2(new_n871), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n873), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n653), .A2(new_n573), .A3(new_n569), .A4(new_n576), .ZN(new_n908));
  INV_X1    g0708(.A(new_n648), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n908), .A2(new_n909), .A3(new_n646), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT26), .B1(new_n653), .B2(new_n634), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n618), .A2(new_n573), .A3(new_n640), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n630), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n679), .B(new_n809), .C1(new_n910), .C2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n807), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n442), .A2(new_n678), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n468), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n442), .B(new_n678), .C1(new_n467), .C2(new_n461), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n914), .A2(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n900), .B1(new_n907), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n899), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n857), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  INV_X1    g0723(.A(new_n809), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n917), .B2(new_n918), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT100), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n729), .A2(new_n733), .ZN(new_n927));
  INV_X1    g0727(.A(new_n720), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT99), .ZN(new_n930));
  INV_X1    g0730(.A(new_n736), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT99), .B1(new_n734), .B2(new_n736), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n929), .A2(new_n678), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n932), .A2(new_n933), .B1(new_n934), .B2(new_n712), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n926), .B1(new_n935), .B2(new_n710), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  AND4_X1   g0737(.A1(new_n926), .A2(new_n937), .A3(new_n710), .A4(new_n735), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n925), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n923), .B1(new_n939), .B2(new_n906), .ZN(new_n940));
  INV_X1    g0740(.A(new_n887), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n869), .A2(new_n870), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n886), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n868), .B1(new_n663), .B2(new_n874), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n892), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n923), .B1(new_n946), .B2(new_n872), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n735), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT100), .B1(new_n948), .B2(new_n711), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n935), .A2(new_n926), .A3(new_n710), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n951), .A3(new_n925), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n537), .A3(new_n951), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(G330), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n953), .B1(new_n537), .B2(new_n951), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n922), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n922), .A2(new_n957), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT101), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n958), .B1(new_n274), .B2(new_n742), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n959), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT101), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n855), .B1(new_n961), .B2(new_n963), .ZN(G367));
  INV_X1    g0764(.A(new_n751), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n758), .B1(new_n206), .B2(new_n416), .C1(new_n228), .C2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n966), .A2(new_n816), .ZN(new_n967));
  INV_X1    g0767(.A(G294), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n781), .A2(new_n968), .B1(new_n783), .B2(new_n790), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n288), .B(new_n969), .C1(G317), .C2(new_n770), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n765), .A2(G116), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT46), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G107), .A2(new_n792), .B1(new_n774), .B2(G303), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT104), .B(G311), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n776), .A2(new_n974), .B1(new_n829), .B2(G97), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n764), .A2(new_n476), .B1(new_n769), .B2(new_n823), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT106), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n288), .B1(new_n762), .B2(new_n378), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(KEYINPUT105), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(KEYINPUT105), .B2(new_n980), .ZN(new_n982));
  INV_X1    g0782(.A(G159), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n781), .A2(new_n983), .B1(new_n783), .B2(new_n233), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G143), .B2(new_n776), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n977), .A2(new_n978), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G68), .A2(new_n792), .B1(new_n774), .B2(G150), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n976), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT47), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n609), .A2(new_n678), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n631), .B(new_n653), .S(new_n991), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n967), .B1(new_n990), .B2(new_n760), .C1(new_n992), .C2(new_n800), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n687), .A2(new_n689), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n689), .A2(new_n685), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n683), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n739), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n567), .A2(new_n568), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n573), .B(new_n569), .C1(new_n1001), .C2(new_n679), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n634), .A2(new_n678), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n690), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT44), .Z(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n690), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n739), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n695), .B(KEYINPUT41), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n746), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1005), .A2(new_n995), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT42), .Z(new_n1019));
  XNOR2_X1  g0819(.A(new_n1004), .B(KEYINPUT102), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n325), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n678), .B1(new_n1022), .B2(new_n573), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1017), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n688), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1020), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1026), .B(new_n1029), .Z(new_n1030));
  OAI21_X1  g0830(.A(new_n993), .B1(new_n1016), .B2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n687), .A2(new_n756), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n693), .A2(new_n206), .A3(new_n288), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(G107), .B2(new_n206), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT107), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n366), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n257), .C1(new_n235), .C2(new_n378), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n751), .B1(new_n225), .B2(new_n257), .C1(new_n693), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1036), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(new_n758), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n764), .A2(new_n378), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n416), .A2(new_n779), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G50), .C2(new_n774), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n783), .A2(new_n235), .B1(new_n769), .B2(new_n368), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n405), .B(new_n1047), .C1(new_n469), .C2(new_n782), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n776), .A2(G159), .B1(new_n829), .B2(G97), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n288), .B1(new_n770), .B2(G326), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n779), .A2(new_n790), .B1(new_n764), .B2(new_n968), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n782), .A2(new_n974), .B1(new_n784), .B2(G303), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n774), .A2(G317), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n789), .C2(new_n777), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT49), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1051), .B1(new_n339), .B2(new_n762), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1050), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n748), .B(new_n1043), .C1(new_n757), .C2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n998), .A2(new_n746), .B1(new_n1032), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n999), .A2(new_n695), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n739), .A2(new_n998), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  XNOR2_X1  g0867(.A(new_n1010), .B(new_n1027), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1013), .B(new_n695), .C1(new_n1068), .C2(new_n1000), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n232), .A2(new_n751), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n758), .C1(new_n331), .C2(new_n206), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n405), .B1(new_n783), .B2(new_n968), .C1(new_n347), .C2(new_n781), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n763), .B(new_n1072), .C1(G116), .C2(new_n792), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n765), .A2(G283), .B1(new_n770), .B2(G322), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT111), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G311), .A2(new_n774), .B1(new_n776), .B2(G317), .ZN(new_n1076));
  XOR2_X1   g0876(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1076), .A2(new_n1077), .B1(KEYINPUT111), .B2(new_n1074), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n1075), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G150), .A2(new_n776), .B1(new_n774), .B2(G159), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT108), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n781), .A2(new_n233), .B1(new_n783), .B2(new_n366), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT109), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n288), .B1(new_n769), .B2(new_n822), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n779), .A2(new_n378), .B1(new_n764), .B2(new_n235), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G87), .C2(new_n829), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1083), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1080), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT112), .Z(new_n1092));
  OAI211_X1 g0892(.A(new_n816), .B(new_n1071), .C1(new_n1092), .C2(new_n760), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1028), .B2(new_n756), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1068), .B2(new_n746), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1069), .A2(new_n1095), .ZN(G390));
  AND3_X1   g0896(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT39), .B1(new_n946), .B2(new_n872), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1097), .A2(new_n1098), .B1(new_n919), .B2(new_n898), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n808), .A2(new_n806), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n704), .A2(new_n679), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n915), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n917), .A2(KEYINPUT113), .A3(new_n918), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT113), .B1(new_n917), .B2(new_n918), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n898), .B1(new_n946), .B2(new_n872), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n917), .A2(new_n918), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n812), .A2(new_n809), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1099), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n925), .B(G330), .C1(new_n936), .C2(new_n938), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT114), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT114), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n951), .A2(new_n1113), .A3(G330), .A4(new_n925), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n807), .B1(new_n706), .B2(new_n809), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1108), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n897), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n895), .A2(new_n1118), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1110), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n746), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n748), .B1(new_n366), .B2(new_n819), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n764), .A2(new_n368), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n781), .A2(new_n823), .B1(new_n783), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n405), .B(new_n1127), .C1(G125), .C2(new_n770), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n774), .A2(G132), .B1(new_n829), .B2(G50), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G159), .A2(new_n792), .B1(new_n776), .B2(G128), .ZN(new_n1130));
  AND4_X1   g0930(.A1(new_n1125), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n781), .A2(new_n297), .B1(new_n783), .B2(new_n331), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1132), .A2(KEYINPUT115), .B1(G283), .B2(new_n776), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(KEYINPUT115), .B2(new_n1132), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT116), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n830), .B1(new_n378), .B2(new_n779), .C1(new_n788), .C2(new_n339), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n405), .B1(new_n769), .B2(new_n968), .C1(new_n837), .C2(new_n764), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1131), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1123), .B1(new_n760), .B2(new_n1139), .C1(new_n896), .C2(new_n755), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1122), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n537), .A2(G330), .A3(new_n951), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n856), .A2(new_n670), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(G330), .B(new_n809), .C1(new_n711), .C2(new_n737), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n915), .B(new_n1101), .C1(new_n1117), .C2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n810), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n951), .A2(new_n1147), .A3(G330), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1117), .A2(new_n1145), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1112), .A2(new_n1114), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1116), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n741), .B1(new_n1156), .B2(new_n1120), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1121), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1141), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(G378));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1143), .B1(new_n1120), .B2(new_n1154), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT120), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1143), .B(KEYINPUT120), .C1(new_n1120), .C2(new_n1154), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n940), .A2(G330), .A3(new_n952), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT119), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n940), .A2(new_n952), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n375), .A2(new_n676), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n404), .B(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1172), .B(new_n1173), .Z(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n1170), .A3(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n953), .A2(KEYINPUT119), .A3(G330), .A4(new_n1174), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n921), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(new_n921), .A3(new_n1177), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1176), .A2(KEYINPUT121), .A3(new_n921), .A4(new_n1177), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1166), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n695), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1174), .A2(new_n754), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n748), .B1(new_n233), .B2(new_n819), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT118), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G150), .A2(new_n792), .B1(new_n776), .B2(G125), .ZN(new_n1194));
  INV_X1    g0994(.A(G128), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n788), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n764), .A2(new_n1126), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n781), .A2(new_n827), .B1(new_n783), .B2(new_n823), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT59), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n829), .A2(G159), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n405), .A2(new_n261), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1044), .A2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT117), .Z(new_n1208));
  AOI22_X1  g1008(.A1(new_n782), .A2(G97), .B1(new_n770), .B2(G283), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n416), .B2(new_n783), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n792), .A2(G68), .B1(new_n829), .B2(G58), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n297), .B2(new_n788), .C1(new_n339), .C2(new_n777), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1206), .B(new_n233), .C1(G33), .C2(G41), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1205), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1193), .B1(new_n1217), .B2(new_n757), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1187), .A2(new_n746), .B1(new_n1191), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1190), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1015), .B(KEYINPUT122), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1156), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT123), .Z(new_n1224));
  INV_X1    g1024(.A(new_n1154), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1149), .A2(new_n754), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n757), .A2(G68), .A3(new_n754), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n777), .A2(new_n968), .B1(new_n764), .B2(new_n331), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G283), .B2(new_n774), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n783), .A2(new_n297), .B1(new_n769), .B2(new_n347), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n288), .B(new_n1230), .C1(G116), .C2(new_n782), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1045), .B1(G77), .B2(new_n829), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n776), .A2(G132), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT125), .Z(new_n1236));
  OAI22_X1  g1036(.A1(new_n781), .A2(new_n1126), .B1(new_n769), .B2(new_n1195), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n405), .B(new_n1237), .C1(G150), .C2(new_n784), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n774), .A2(G137), .B1(new_n829), .B2(G58), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n792), .A2(G50), .B1(new_n765), .B2(G159), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1234), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n748), .B(new_n1227), .C1(new_n1243), .C2(new_n757), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1225), .A2(new_n746), .B1(new_n1226), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1224), .A2(new_n1245), .ZN(G381));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G387), .A2(new_n1249), .A3(G378), .A4(new_n1250), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n1251), .A2(G375), .A3(G381), .ZN(G407));
  INV_X1    g1052(.A(G213), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G343), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1159), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G375), .C2(new_n1255), .ZN(G409));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(new_n1247), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G387), .A2(new_n1247), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1261), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1219), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1183), .A2(new_n746), .A3(new_n1184), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1187), .A2(new_n1188), .A3(new_n1222), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1191), .A2(new_n1218), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1159), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1254), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1221), .B1(new_n1155), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n1154), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n695), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(G384), .A3(new_n1245), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1277), .B2(new_n1245), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT62), .B1(new_n1273), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1254), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1286), .B(new_n1254), .C1(new_n1267), .C2(new_n1272), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1281), .A2(KEYINPUT62), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1282), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1280), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1291), .A2(new_n1278), .B1(G2897), .B2(new_n1254), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1254), .A2(G2897), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1279), .A2(new_n1280), .A3(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1266), .B1(new_n1290), .B2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1265), .B(new_n1298), .C1(new_n1273), .C2(new_n1295), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT63), .B1(new_n1273), .B2(new_n1281), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1281), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1300), .A2(new_n1305), .ZN(G405));
  AOI21_X1  g1106(.A(G378), .B1(new_n1190), .B2(new_n1219), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1267), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1281), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1281), .A2(new_n1310), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT127), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1312), .B(new_n1313), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(new_n1265), .ZN(G402));
endmodule


