

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592;

  OR2_X1 U322 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U323 ( .A(G43GAT), .B(G190GAT), .ZN(n318) );
  XNOR2_X1 U324 ( .A(n318), .B(G134GAT), .ZN(n444) );
  XNOR2_X1 U325 ( .A(G36GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U326 ( .A(n319), .B(KEYINPUT75), .ZN(n410) );
  XNOR2_X1 U327 ( .A(n553), .B(KEYINPUT36), .ZN(n504) );
  XOR2_X2 U328 ( .A(n334), .B(n333), .Z(n571) );
  XNOR2_X1 U329 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U330 ( .A(KEYINPUT64), .B(n424), .Z(n290) );
  XOR2_X1 U331 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n291) );
  XOR2_X1 U332 ( .A(n463), .B(n462), .Z(n292) );
  XNOR2_X1 U333 ( .A(n355), .B(n354), .ZN(n356) );
  INV_X1 U334 ( .A(n561), .ZN(n393) );
  INV_X1 U335 ( .A(KEYINPUT33), .ZN(n364) );
  AND2_X1 U336 ( .A1(n394), .A2(n393), .ZN(n401) );
  XNOR2_X1 U337 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U338 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U339 ( .A(n581), .B(KEYINPUT41), .ZN(n563) );
  XOR2_X1 U340 ( .A(n371), .B(n370), .Z(n581) );
  XOR2_X1 U341 ( .A(n392), .B(n391), .Z(n561) );
  XNOR2_X1 U342 ( .A(n467), .B(G190GAT), .ZN(n468) );
  XNOR2_X1 U343 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n294) );
  XNOR2_X1 U345 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n313) );
  XOR2_X1 U347 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n296) );
  XNOR2_X1 U348 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U350 ( .A(G155GAT), .B(G148GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(G120GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n311) );
  XOR2_X1 U354 ( .A(G113GAT), .B(KEYINPUT0), .Z(n452) );
  XOR2_X1 U355 ( .A(G85GAT), .B(G162GAT), .Z(n302) );
  XNOR2_X1 U356 ( .A(G29GAT), .B(G134GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U358 ( .A(n452), .B(n303), .Z(n305) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U361 ( .A(n306), .B(G57GAT), .Z(n309) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n307), .B(KEYINPUT2), .ZN(n427) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(n427), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U367 ( .A(n313), .B(n312), .Z(n473) );
  INV_X1 U368 ( .A(n473), .ZN(n529) );
  XOR2_X1 U369 ( .A(G92GAT), .B(G85GAT), .Z(n315) );
  XNOR2_X1 U370 ( .A(G99GAT), .B(G106GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n363) );
  XNOR2_X1 U372 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n316) );
  XOR2_X1 U373 ( .A(n316), .B(KEYINPUT8), .Z(n374) );
  INV_X1 U374 ( .A(n374), .ZN(n317) );
  XOR2_X1 U375 ( .A(n363), .B(n317), .Z(n334) );
  XNOR2_X1 U376 ( .A(n444), .B(n410), .ZN(n325) );
  XOR2_X1 U377 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n321) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n323) );
  INV_X1 U380 ( .A(KEYINPUT9), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n327) );
  INV_X1 U383 ( .A(KEYINPUT76), .ZN(n326) );
  NAND2_X1 U384 ( .A1(n327), .A2(n326), .ZN(n330) );
  INV_X1 U385 ( .A(n327), .ZN(n328) );
  NAND2_X1 U386 ( .A1(n328), .A2(KEYINPUT76), .ZN(n329) );
  NAND2_X1 U387 ( .A1(n330), .A2(n329), .ZN(n332) );
  XOR2_X1 U388 ( .A(G50GAT), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U389 ( .A(n433), .B(KEYINPUT74), .ZN(n331) );
  XOR2_X2 U390 ( .A(KEYINPUT77), .B(n571), .Z(n553) );
  XOR2_X1 U391 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n336) );
  XNOR2_X1 U392 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n353) );
  XOR2_X1 U394 ( .A(G211GAT), .B(G78GAT), .Z(n338) );
  XNOR2_X1 U395 ( .A(G183GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n340) );
  XNOR2_X1 U398 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U400 ( .A(n342), .B(n341), .Z(n347) );
  XOR2_X1 U401 ( .A(G1GAT), .B(G8GAT), .Z(n386) );
  XOR2_X1 U402 ( .A(G22GAT), .B(G155GAT), .Z(n432) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .Z(n447) );
  XOR2_X1 U404 ( .A(n432), .B(n447), .Z(n344) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n386), .B(n345), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U409 ( .A(n348), .B(KEYINPUT12), .Z(n351) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n291), .B(n349), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n360), .B(KEYINPUT79), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n587) );
  INV_X1 U415 ( .A(n587), .ZN(n568) );
  NAND2_X1 U416 ( .A1(n504), .A2(n568), .ZN(n357) );
  XOR2_X1 U417 ( .A(KEYINPUT45), .B(KEYINPUT107), .Z(n355) );
  INV_X1 U418 ( .A(KEYINPUT65), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n372) );
  XOR2_X1 U420 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n359) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(KEYINPUT72), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n371) );
  XOR2_X1 U423 ( .A(G148GAT), .B(G78GAT), .Z(n436) );
  XOR2_X1 U424 ( .A(G204GAT), .B(G64GAT), .Z(n414) );
  XNOR2_X1 U425 ( .A(n436), .B(n414), .ZN(n369) );
  XOR2_X1 U426 ( .A(G120GAT), .B(G71GAT), .Z(n451) );
  XOR2_X1 U427 ( .A(n451), .B(n360), .Z(n362) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n363), .B(KEYINPUT73), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  INV_X1 U432 ( .A(n581), .ZN(n472) );
  NOR2_X1 U433 ( .A1(n372), .A2(n472), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n373), .B(KEYINPUT108), .ZN(n394) );
  XNOR2_X1 U435 ( .A(n374), .B(KEYINPUT68), .ZN(n376) );
  NAND2_X1 U436 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n392) );
  XOR2_X1 U438 ( .A(KEYINPUT67), .B(G197GAT), .Z(n378) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(G141GAT), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n380) );
  XNOR2_X1 U442 ( .A(KEYINPUT66), .B(KEYINPUT69), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n390) );
  XOR2_X1 U445 ( .A(G113GAT), .B(G43GAT), .Z(n384) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(G50GAT), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U448 ( .A(n385), .B(G15GAT), .Z(n388) );
  XNOR2_X1 U449 ( .A(G169GAT), .B(n386), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n563), .A2(n561), .ZN(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT46), .B(KEYINPUT106), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U455 ( .A1(n397), .A2(n587), .ZN(n398) );
  NOR2_X1 U456 ( .A1(n571), .A2(n398), .ZN(n399) );
  XOR2_X1 U457 ( .A(KEYINPUT47), .B(n399), .Z(n400) );
  XNOR2_X2 U458 ( .A(n402), .B(KEYINPUT48), .ZN(n558) );
  XOR2_X1 U459 ( .A(G176GAT), .B(G183GAT), .Z(n404) );
  XNOR2_X1 U460 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT17), .B(KEYINPUT87), .Z(n406) );
  XNOR2_X1 U463 ( .A(KEYINPUT86), .B(KEYINPUT18), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U465 ( .A(n408), .B(n407), .Z(n456) );
  INV_X1 U466 ( .A(n456), .ZN(n420) );
  XNOR2_X1 U467 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n409), .B(G211GAT), .ZN(n434) );
  XNOR2_X1 U469 ( .A(n410), .B(n434), .ZN(n418) );
  XOR2_X1 U470 ( .A(KEYINPUT94), .B(G92GAT), .Z(n412) );
  XNOR2_X1 U471 ( .A(G8GAT), .B(G190GAT), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U473 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n479) );
  NAND2_X1 U478 ( .A1(n558), .A2(n479), .ZN(n422) );
  XOR2_X1 U479 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  NAND2_X1 U481 ( .A1(n529), .A2(n423), .ZN(n424) );
  XOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n426) );
  XNOR2_X1 U483 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U485 ( .A(n427), .B(G204GAT), .Z(n429) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n441) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U491 ( .A(n437), .B(n436), .Z(n439) );
  XNOR2_X1 U492 ( .A(G218GAT), .B(G106GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n482) );
  NAND2_X1 U495 ( .A1(n290), .A2(n482), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n457) );
  XOR2_X1 U498 ( .A(n444), .B(KEYINPUT85), .Z(n446) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U501 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U503 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U506 ( .A(n456), .B(n455), .Z(n480) );
  NAND2_X1 U507 ( .A1(n457), .A2(n480), .ZN(n465) );
  NOR2_X1 U508 ( .A1(n465), .A2(n587), .ZN(n459) );
  INV_X1 U509 ( .A(G183GAT), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  NOR2_X1 U511 ( .A1(n393), .A2(n465), .ZN(n461) );
  INV_X1 U512 ( .A(G169GAT), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n461), .B(n460), .ZN(G1348GAT) );
  INV_X1 U514 ( .A(n563), .ZN(n518) );
  NOR2_X1 U515 ( .A1(n465), .A2(n518), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n463) );
  XNOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n464), .B(n292), .ZN(G1349GAT) );
  INV_X1 U519 ( .A(n465), .ZN(n466) );
  NAND2_X1 U520 ( .A1(n466), .A2(n553), .ZN(n469) );
  XOR2_X1 U521 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n467) );
  XOR2_X1 U522 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n471) );
  XNOR2_X1 U523 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n470) );
  XNOR2_X1 U524 ( .A(n471), .B(n470), .ZN(n494) );
  NOR2_X1 U525 ( .A1(n393), .A2(n472), .ZN(n507) );
  XNOR2_X1 U526 ( .A(n482), .B(KEYINPUT28), .ZN(n537) );
  INV_X1 U527 ( .A(n537), .ZN(n474) );
  INV_X1 U528 ( .A(n479), .ZN(n532) );
  XOR2_X1 U529 ( .A(KEYINPUT27), .B(n532), .Z(n478) );
  NAND2_X1 U530 ( .A1(n473), .A2(n478), .ZN(n560) );
  NOR2_X1 U531 ( .A1(n474), .A2(n560), .ZN(n540) );
  INV_X1 U532 ( .A(n480), .ZN(n542) );
  XNOR2_X1 U533 ( .A(n542), .B(KEYINPUT88), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n540), .A2(n475), .ZN(n488) );
  NOR2_X1 U535 ( .A1(n480), .A2(n482), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT95), .B(n476), .Z(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT26), .B(n477), .ZN(n575) );
  NAND2_X1 U538 ( .A1(n575), .A2(n478), .ZN(n485) );
  NAND2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT25), .B(n483), .Z(n484) );
  NAND2_X1 U542 ( .A1(n485), .A2(n484), .ZN(n486) );
  NAND2_X1 U543 ( .A1(n486), .A2(n529), .ZN(n487) );
  NAND2_X1 U544 ( .A1(n488), .A2(n487), .ZN(n502) );
  NOR2_X1 U545 ( .A1(n553), .A2(n587), .ZN(n490) );
  XNOR2_X1 U546 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U548 ( .A1(n502), .A2(n491), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT96), .B(n492), .Z(n519) );
  NAND2_X1 U550 ( .A1(n507), .A2(n519), .ZN(n500) );
  NOR2_X1 U551 ( .A1(n529), .A2(n500), .ZN(n493) );
  XOR2_X1 U552 ( .A(n494), .B(n493), .Z(G1324GAT) );
  NOR2_X1 U553 ( .A1(n532), .A2(n500), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U556 ( .A1(n542), .A2(n500), .ZN(n498) );
  XNOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U560 ( .A1(n537), .A2(n500), .ZN(n501) );
  XOR2_X1 U561 ( .A(G22GAT), .B(n501), .Z(G1327GAT) );
  NAND2_X1 U562 ( .A1(n587), .A2(n502), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n503), .B(KEYINPUT101), .ZN(n505) );
  NAND2_X1 U564 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(KEYINPUT37), .B(n506), .ZN(n528) );
  NAND2_X1 U566 ( .A1(n507), .A2(n528), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n508), .B(KEYINPUT38), .ZN(n516) );
  NOR2_X1 U568 ( .A1(n516), .A2(n529), .ZN(n510) );
  XNOR2_X1 U569 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(n511), .ZN(G1328GAT) );
  XNOR2_X1 U572 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n513) );
  NOR2_X1 U573 ( .A1(n532), .A2(n516), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n513), .B(n512), .ZN(G1329GAT) );
  NOR2_X1 U575 ( .A1(n516), .A2(n542), .ZN(n514) );
  XOR2_X1 U576 ( .A(n514), .B(KEYINPUT40), .Z(n515) );
  XNOR2_X1 U577 ( .A(G43GAT), .B(n515), .ZN(G1330GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n537), .ZN(n517) );
  XOR2_X1 U579 ( .A(G50GAT), .B(n517), .Z(G1331GAT) );
  NOR2_X1 U580 ( .A1(n561), .A2(n518), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n527), .A2(n519), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n529), .A2(n524), .ZN(n520) );
  XOR2_X1 U583 ( .A(G57GAT), .B(n520), .Z(n521) );
  XNOR2_X1 U584 ( .A(KEYINPUT42), .B(n521), .ZN(G1332GAT) );
  NOR2_X1 U585 ( .A1(n532), .A2(n524), .ZN(n522) );
  XOR2_X1 U586 ( .A(G64GAT), .B(n522), .Z(G1333GAT) );
  NOR2_X1 U587 ( .A1(n542), .A2(n524), .ZN(n523) );
  XOR2_X1 U588 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U589 ( .A1(n537), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n529), .A2(n536), .ZN(n530) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n530), .Z(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT104), .B(n531), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n536), .ZN(n534) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(KEYINPUT105), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n542), .A2(n536), .ZN(n535) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  XOR2_X1 U604 ( .A(G113GAT), .B(KEYINPUT109), .Z(n544) );
  NAND2_X1 U605 ( .A1(n558), .A2(n540), .ZN(n541) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n554), .A2(n561), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n546) );
  NAND2_X1 U610 ( .A1(n554), .A2(n563), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT110), .Z(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n568), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G134GAT), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n575), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n572) );
  NAND2_X1 U625 ( .A1(n572), .A2(n561), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n565) );
  NAND2_X1 U628 ( .A1(n572), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT52), .Z(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n572), .A2(n568), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(KEYINPUT116), .ZN(n570) );
  XNOR2_X1 U634 ( .A(G155GAT), .B(n570), .ZN(G1346GAT) );
  XOR2_X1 U635 ( .A(G162GAT), .B(KEYINPUT117), .Z(n574) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n574), .B(n573), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n290), .A2(n575), .ZN(n589) );
  NOR2_X1 U639 ( .A1(n393), .A2(n589), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n577) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT122), .B(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n589), .ZN(n586) );
  XOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT124), .B(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n589), .ZN(n588) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
  INV_X1 U653 ( .A(n589), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n504), .A2(n590), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

