//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT92), .B1(new_n209), .B2(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(G43gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n210), .B(new_n213), .C1(G43gat), .C2(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT93), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT94), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n209), .A2(G50gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n212), .A2(G43gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT90), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n225), .B2(new_n226), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(KEYINPUT15), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G29gat), .A2(G36gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n224), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n222), .A2(KEYINPUT91), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n222), .A2(KEYINPUT91), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n221), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n236), .A2(new_n232), .ZN(new_n237));
  OAI22_X1  g036(.A1(new_n217), .A2(new_n233), .B1(new_n237), .B2(new_n231), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT96), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n231), .B1(new_n232), .B2(new_n236), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n224), .A2(new_n231), .A3(new_n232), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT93), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n216), .B(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n241), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT96), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT17), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G15gat), .B(G22gat), .ZN(new_n249));
  INV_X1    g048(.A(G1gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT16), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252));
  OAI221_X1 g051(.A(new_n251), .B1(new_n252), .B2(G8gat), .C1(new_n250), .C2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(G8gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(new_n238), .B2(new_n239), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT97), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(KEYINPUT18), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G229gat), .A2(G233gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n255), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n257), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n253), .B(new_n254), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n245), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n262), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n261), .B(KEYINPUT13), .Z(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n248), .A2(new_n256), .B1(new_n238), .B2(new_n255), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n260), .B1(new_n270), .B2(new_n261), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n208), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n261), .A3(new_n262), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n259), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n274), .A2(new_n268), .A3(new_n263), .A4(new_n207), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277));
  XOR2_X1   g076(.A(G1gat), .B(G29gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT0), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT2), .B1(new_n287), .B2(KEYINPUT76), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n286), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n287), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n282), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(new_n295), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT76), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(new_n294), .A3(new_n297), .ZN(new_n308));
  OR3_X1    g107(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n309), .A2(new_n283), .B1(G155gat), .B2(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n302), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n315));
  OAI21_X1  g114(.A(G134gat), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(G127gat), .A2(G134gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n317), .C1(KEYINPUT1), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G120gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT66), .ZN(new_n324));
  OR3_X1    g123(.A1(new_n322), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n304), .A2(new_n313), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n311), .A2(new_n302), .A3(new_n328), .A4(new_n319), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n334));
  AND2_X1   g133(.A1(new_n319), .A2(new_n328), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n308), .A2(new_n310), .B1(new_n296), .B2(new_n301), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n330), .B(new_n331), .C1(new_n333), .C2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n339));
  NAND2_X1  g138(.A1(new_n311), .A2(new_n302), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n329), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n332), .ZN(new_n342));
  INV_X1    g141(.A(new_n331), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n334), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n335), .A2(new_n336), .A3(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n347), .A2(new_n339), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n335), .B1(new_n340), .B2(KEYINPUT3), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n343), .B1(new_n351), .B2(new_n313), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n281), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n277), .B1(new_n354), .B2(KEYINPUT6), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n338), .A2(new_n344), .B1(new_n350), .B2(new_n352), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n357));
  NOR4_X1   g156(.A1(new_n356), .A2(KEYINPUT85), .A3(new_n357), .A4(new_n281), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT72), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(KEYINPUT72), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n368), .A2(new_n360), .A3(new_n364), .A4(new_n362), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT73), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT73), .B1(new_n367), .B2(new_n369), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G226gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT26), .ZN(new_n377));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n376), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G183gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT27), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G183gat), .ZN(new_n388));
  INV_X1    g187(.A(G190gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT27), .B(G183gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT28), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n384), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n376), .A2(KEYINPUT23), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n396), .A2(new_n380), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n378), .ZN(new_n401));
  NAND3_X1  g200(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT25), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n396), .A2(KEYINPUT25), .A3(new_n398), .A4(new_n380), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n406), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n400), .A2(new_n378), .B1(new_n402), .B2(KEYINPUT64), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n395), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n375), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n402), .A2(KEYINPUT64), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n401), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT25), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n380), .A3(new_n398), .ZN(new_n417));
  AND2_X1   g216(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n378), .A2(new_n400), .B1(new_n418), .B2(G190gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n391), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n393), .A2(KEYINPUT28), .A3(new_n389), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n415), .A2(new_n420), .B1(new_n423), .B2(new_n384), .ZN(new_n424));
  INV_X1    g223(.A(new_n375), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n372), .B1(new_n412), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n424), .B2(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n375), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n367), .A2(new_n369), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT73), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(new_n428), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT38), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n412), .A2(new_n372), .A3(new_n426), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n435), .B1(new_n429), .B2(new_n430), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT37), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n444), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n442), .A2(new_n445), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n345), .A2(new_n353), .ZN(new_n448));
  INV_X1    g247(.A(new_n281), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT6), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n356), .A2(new_n281), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT84), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n357), .B1(new_n356), .B2(new_n281), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n345), .A2(new_n353), .A3(new_n281), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n359), .B(new_n447), .C1(new_n452), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT86), .ZN(new_n458));
  INV_X1    g257(.A(new_n354), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n459), .A2(KEYINPUT84), .A3(new_n451), .A4(new_n357), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n359), .A4(new_n447), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT74), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n443), .B2(new_n444), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n427), .A2(KEYINPUT74), .A3(new_n436), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT37), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  INV_X1    g268(.A(new_n440), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n437), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT38), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n464), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n330), .A2(new_n349), .A3(new_n347), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(KEYINPUT83), .A3(new_n343), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT83), .B1(new_n477), .B2(new_n343), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n342), .A2(new_n343), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n476), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n485), .A3(new_n281), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n427), .A2(new_n440), .A3(new_n436), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n446), .A2(KEYINPUT30), .A3(new_n440), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT40), .A4(new_n281), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n488), .A2(new_n459), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT29), .B1(new_n336), .B2(new_n312), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT80), .B1(new_n435), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n313), .A2(new_n411), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n372), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT29), .B1(new_n367), .B2(new_n369), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n340), .B1(new_n503), .B2(KEYINPUT3), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT79), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT79), .B(new_n340), .C1(new_n503), .C2(KEYINPUT3), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n499), .A2(new_n502), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n509), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(new_n504), .C1(new_n435), .C2(new_n498), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT81), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n372), .A2(new_n501), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT81), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n512), .A4(new_n504), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n510), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n511), .B1(new_n510), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n497), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n510), .A2(new_n518), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G22gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n510), .A2(new_n511), .A3(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT82), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G78gat), .B(G106gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G50gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(KEYINPUT82), .A3(new_n524), .A4(new_n528), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n496), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n475), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n354), .A2(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n450), .A2(new_n451), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n494), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n415), .A2(new_n420), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n335), .A3(new_n395), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT68), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n424), .A2(new_n543), .A3(new_n335), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n410), .A2(new_n329), .ZN(new_n545));
  NAND2_X1  g344(.A1(G227gat), .A2(G233gat), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT34), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n551));
  INV_X1    g350(.A(new_n546), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT33), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT69), .B(G71gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G99gat), .ZN(new_n556));
  XOR2_X1   g355(.A(G15gat), .B(G43gat), .Z(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  AOI221_X4 g359(.A(new_n550), .B1(KEYINPUT33), .B2(new_n558), .C1(new_n551), .C2(new_n552), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n549), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n551), .A2(new_n552), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n553), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n561), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n548), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n563), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT71), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n548), .A2(KEYINPUT70), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n562), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n562), .B2(new_n570), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT36), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n533), .A2(new_n539), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n530), .A2(new_n531), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n570), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n462), .A2(new_n359), .ZN(new_n584));
  INV_X1    g383(.A(new_n494), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT88), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n587));
  AOI211_X1 g386(.A(new_n587), .B(new_n494), .C1(new_n462), .C2(new_n359), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n580), .B(new_n583), .C1(new_n586), .C2(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n530), .B(new_n531), .C1(new_n575), .C2(new_n576), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT35), .B1(new_n590), .B2(new_n538), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n276), .B1(new_n579), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT102), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT7), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT103), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n602), .A2(new_n604), .A3(G85gat), .A4(G92gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT8), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(KEYINPUT103), .A3(new_n603), .ZN(new_n609));
  OR2_X1    g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n605), .A2(new_n607), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n248), .B(new_n613), .C1(KEYINPUT17), .C2(new_n245), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n238), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G190gat), .B(G218gat), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n600), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n617), .A2(new_n618), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n598), .B(new_n599), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G71gat), .B(G78gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT9), .ZN(new_n630));
  INV_X1    g429(.A(G71gat), .ZN(new_n631));
  INV_X1    g430(.A(G78gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G57gat), .ZN(new_n634));
  INV_X1    g433(.A(G64gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G57gat), .A2(G64gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n627), .A2(new_n628), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(KEYINPUT99), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n642));
  OAI21_X1  g441(.A(G64gat), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n635), .B1(new_n644), .B2(new_n634), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n643), .A2(new_n633), .A3(new_n627), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(KEYINPUT21), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n264), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT101), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT21), .B1(new_n640), .B2(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G127gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G155gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n654), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n640), .A2(new_n646), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n613), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n611), .A2(new_n612), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n611), .A2(new_n612), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n640), .A3(new_n646), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n613), .A2(new_n665), .A3(new_n663), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n662), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT105), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n664), .A2(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n662), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n675), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n661), .B(KEYINPUT106), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n677), .ZN(new_n685));
  INV_X1    g484(.A(new_n680), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n626), .A2(new_n660), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n593), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n536), .A2(new_n535), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G8gat), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n691), .A2(new_n494), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(G8gat), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n691), .B2(new_n494), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT42), .B2(new_n698), .ZN(G1325gat));
  INV_X1    g501(.A(new_n691), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n703), .B2(new_n578), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n582), .A2(G15gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(G1326gat));
  NOR2_X1   g505(.A1(new_n593), .A2(new_n580), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n622), .A2(new_n625), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n659), .A3(new_n688), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT108), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n712), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n593), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n659), .A2(new_n689), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n626), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(new_n219), .A3(new_n693), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n475), .A2(new_n532), .B1(new_n573), .B2(new_n577), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n534), .B2(new_n538), .ZN(new_n725));
  AOI211_X1 g524(.A(KEYINPUT109), .B(new_n537), .C1(new_n530), .C2(new_n531), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n723), .A2(new_n727), .B1(new_n591), .B2(new_n589), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n722), .B1(new_n728), .B2(new_n626), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n626), .A2(new_n722), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n579), .B2(new_n592), .ZN(new_n731));
  INV_X1    g530(.A(new_n276), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n718), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n692), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n721), .A2(new_n735), .ZN(G1328gat));
  NAND4_X1  g535(.A1(new_n717), .A2(new_n220), .A3(new_n494), .A4(new_n719), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT46), .Z(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n734), .B2(new_n585), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  NAND3_X1  g539(.A1(new_n717), .A2(new_n581), .A3(new_n719), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n209), .ZN(new_n742));
  INV_X1    g541(.A(new_n578), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n734), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g545(.A(G50gat), .B1(new_n734), .B2(new_n580), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n718), .A2(new_n626), .A3(G50gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n707), .A2(new_n748), .B1(KEYINPUT110), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1331gat));
  NAND3_X1  g552(.A1(new_n626), .A2(new_n660), .A3(new_n688), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n728), .A2(new_n276), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n693), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT99), .B(G57gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1332gat));
  XOR2_X1   g557(.A(new_n494), .B(KEYINPUT111), .Z(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n765), .B(new_n767), .ZN(G1333gat));
  NAND3_X1  g567(.A1(new_n755), .A2(new_n631), .A3(new_n581), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n755), .A2(new_n743), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n631), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n534), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n732), .A2(new_n659), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT114), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n723), .A2(new_n727), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n708), .B(new_n776), .C1(new_n777), .C2(new_n592), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n728), .A2(new_n626), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n776), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n779), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n689), .A2(G85gat), .A3(new_n692), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n776), .A2(new_n688), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n729), .A2(new_n731), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n692), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1336gat));
  NOR3_X1   g590(.A1(new_n759), .A2(G92gat), .A3(new_n689), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n784), .A2(new_n785), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  OAI21_X1  g593(.A(G92gat), .B1(new_n789), .B2(new_n759), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n789), .A2(new_n585), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n797), .A2(G92gat), .B1(new_n798), .B2(new_n792), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(new_n794), .ZN(G1337gat));
  NOR3_X1   g599(.A1(new_n582), .A2(G99gat), .A3(new_n689), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G99gat), .B1(new_n789), .B2(new_n578), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1338gat));
  NOR3_X1   g603(.A1(new_n580), .A2(G106gat), .A3(new_n689), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n785), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n729), .A2(new_n534), .A3(new_n731), .A4(new_n788), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT53), .B1(new_n807), .B2(G106gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n807), .A2(new_n810), .A3(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n807), .B2(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n805), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n780), .B2(new_n782), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n809), .B1(new_n815), .B2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n671), .B2(new_n683), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n674), .B2(new_n673), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n671), .A2(new_n821), .A3(new_n683), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n686), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n818), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n822), .A2(new_n686), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n671), .A2(new_n672), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(new_n661), .A3(new_n674), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n825), .B(KEYINPUT55), .C1(new_n827), .C2(new_n819), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n824), .A2(new_n828), .A3(new_n681), .ZN(new_n829));
  INV_X1    g628(.A(new_n206), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n270), .A2(new_n261), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n266), .A2(new_n267), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n275), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n708), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n834), .A2(new_n688), .B1(new_n276), .B2(new_n829), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n708), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n659), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n709), .A2(new_n732), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n590), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n693), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n759), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n322), .A3(new_n276), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n692), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n840), .A2(new_n580), .A3(new_n581), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n732), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n850), .B2(new_n851), .ZN(G1340gat));
  NOR3_X1   g651(.A1(new_n847), .A2(new_n320), .A3(new_n689), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n844), .A2(new_n688), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n320), .ZN(G1341gat));
  NOR3_X1   g654(.A1(new_n659), .A2(new_n315), .A3(new_n314), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n844), .A2(new_n856), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n847), .A2(new_n659), .B1(new_n315), .B2(new_n314), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1342gat));
  NAND2_X1  g658(.A1(new_n708), .A2(new_n585), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT118), .Z(new_n861));
  OR3_X1    g660(.A1(new_n842), .A2(G134gat), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n847), .B2(new_n626), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  NAND3_X1  g665(.A1(new_n824), .A2(new_n828), .A3(new_n681), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n272), .B2(new_n275), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n275), .A2(new_n688), .A3(new_n833), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n276), .A2(new_n829), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n869), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n874), .A3(new_n626), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n660), .B1(new_n875), .B2(new_n835), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n690), .A2(new_n276), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n534), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n626), .B1(new_n868), .B2(new_n870), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n660), .B1(new_n881), .B2(new_n835), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n534), .C1(new_n882), .C2(new_n877), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n578), .A2(new_n846), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n732), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n743), .A2(new_n580), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n840), .A2(new_n693), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n276), .A2(new_n289), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT121), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n889), .A2(new_n843), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n887), .B(new_n892), .C1(KEYINPUT120), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n892), .B2(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n883), .A2(new_n884), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(KEYINPUT57), .B2(new_n878), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n289), .B1(new_n897), .B2(new_n276), .ZN(new_n898));
  INV_X1    g697(.A(new_n892), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n894), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(new_n889), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n902), .A2(new_n290), .A3(new_n688), .A4(new_n759), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n290), .C1(new_n897), .C2(new_n688), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n708), .B1(new_n836), .B2(new_n873), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n626), .A2(new_n867), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n907), .A2(new_n871), .B1(new_n834), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n906), .B(new_n839), .C1(new_n909), .C2(new_n660), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n876), .B2(new_n877), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n580), .A2(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n840), .A2(new_n534), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n913), .A2(new_n688), .A3(new_n915), .A4(new_n884), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n905), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n903), .B1(new_n904), .B2(new_n917), .ZN(G1345gat));
  NOR2_X1   g717(.A1(new_n659), .A2(new_n298), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n897), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n660), .A3(new_n759), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n298), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n921), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1346gat));
  AOI21_X1  g727(.A(new_n299), .B1(new_n897), .B2(new_n708), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n889), .A2(G162gat), .A3(new_n861), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G162gat), .B1(new_n886), .B2(new_n626), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  INV_X1    g732(.A(new_n930), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n693), .A2(new_n585), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n840), .A2(new_n580), .A3(new_n581), .A4(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G169gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(new_n732), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n693), .B1(new_n838), .B2(new_n839), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n590), .A2(new_n759), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n276), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n940), .B1(new_n939), .B2(new_n945), .ZN(G1348gat));
  OAI21_X1  g745(.A(G176gat), .B1(new_n938), .B2(new_n689), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n689), .A2(G176gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n943), .B2(new_n948), .ZN(G1349gat));
  AND2_X1   g748(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n950));
  OAI21_X1  g749(.A(G183gat), .B1(new_n938), .B2(new_n659), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n941), .A2(new_n393), .A3(new_n660), .A4(new_n942), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT127), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n944), .A2(new_n389), .A3(new_n708), .ZN(new_n957));
  OAI21_X1  g756(.A(G190gat), .B1(new_n938), .B2(new_n626), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1351gat));
  AND3_X1   g761(.A1(new_n941), .A2(new_n843), .A3(new_n888), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n276), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n913), .A2(new_n915), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n578), .A2(new_n937), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n276), .A2(G197gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n688), .A3(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G204gat), .ZN(new_n971));
  INV_X1    g770(.A(G204gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n963), .A2(new_n972), .A3(new_n688), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n975), .ZN(G1353gat));
  INV_X1    g775(.A(G211gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n963), .A2(new_n977), .A3(new_n660), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n913), .A2(new_n660), .A3(new_n915), .A4(new_n966), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n708), .A3(new_n966), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G218gat), .ZN(new_n984));
  INV_X1    g783(.A(G218gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n963), .A2(new_n985), .A3(new_n708), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1355gat));
endmodule


