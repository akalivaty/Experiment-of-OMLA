//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n440, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(new_n440), .A2(G57), .A3(G69), .A4(G108), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2106), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT70), .B1(new_n471), .B2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(G137), .A3(new_n469), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(G2104), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n470), .A2(new_n477), .A3(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n476), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n476), .A2(new_n469), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n474), .A2(G126), .A3(G2105), .A4(new_n475), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n474), .A2(G138), .A3(new_n469), .A4(new_n475), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT3), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n473), .A3(new_n501), .A4(new_n469), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n467), .A2(new_n504), .A3(new_n469), .A4(new_n499), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI211_X1 g081(.A(KEYINPUT73), .B(new_n495), .C1(new_n497), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n509));
  INV_X1    g084(.A(new_n495), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT75), .A3(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(new_n518), .B1(KEYINPUT5), .B2(new_n515), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n523), .B1(new_n521), .B2(KEYINPUT74), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT6), .A3(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n515), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n526), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(G88), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n522), .A2(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(new_n519), .A2(new_n529), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n527), .A2(G51), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n535), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AOI22_X1  g116(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n527), .A2(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n530), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n527), .A2(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n530), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n519), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n521), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT77), .Z(G176));
  XOR2_X1   g133(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n564));
  INV_X1    g139(.A(new_n518), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT75), .B1(new_n517), .B2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n534), .A2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n527), .A2(G53), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  XNOR2_X1  g152(.A(G171), .B(new_n577), .ZN(G301));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n534), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n527), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n519), .A2(G86), .A3(new_n529), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n527), .A2(G48), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n521), .ZN(G305));
  AOI22_X1  g162(.A1(new_n534), .A2(G85), .B1(G47), .B2(new_n527), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n567), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n530), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n595), .A2(new_n598), .B1(G54), .B2(new_n527), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n567), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(G868), .B2(new_n606), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT81), .ZN(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(new_n575), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n572), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n606), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n479), .A2(new_n467), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n483), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n486), .A2(G135), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n623), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n636), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT17), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n666));
  INV_X1    g241(.A(new_n661), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  AOI22_X1  g243(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n661), .A3(new_n664), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n669), .B(new_n671), .C1(new_n665), .C2(new_n666), .ZN(new_n672));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G23), .ZN(new_n680));
  AND3_X1   g255(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT33), .Z(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT87), .B(G16), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G1971), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n679), .A2(G6), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n584), .A2(new_n585), .ZN(new_n690));
  OAI211_X1 g265(.A(G61), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n691));
  NAND2_X1  g266(.A1(G73), .A2(G543), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n521), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n689), .B1(new_n694), .B2(new_n679), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n697), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n698), .B(new_n699), .C1(new_n687), .C2(G1971), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n683), .B2(G1976), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n684), .A2(new_n688), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT89), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT89), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(KEYINPUT34), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n486), .A2(G131), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT86), .ZN(new_n709));
  OR2_X1    g284(.A1(G95), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n483), .A2(G119), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n707), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n705), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n703), .A2(new_n704), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(new_n685), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT88), .B(G1986), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n719), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n719), .A2(new_n728), .A3(new_n722), .A4(new_n725), .ZN(new_n732));
  INV_X1    g307(.A(new_n685), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n554), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT91), .B(G1341), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n486), .A2(G139), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT93), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(new_n469), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AND3_X1   g318(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G33), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n706), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n706), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT29), .Z(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n606), .A2(new_n679), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G4), .B2(new_n679), .ZN(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n750), .A2(new_n751), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  NOR2_X1   g337(.A1(G27), .A2(G29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G164), .B2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G2078), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n679), .A2(G5), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G171), .B2(new_n679), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT97), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n733), .A2(KEYINPUT23), .A3(G20), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT23), .ZN(new_n772));
  INV_X1    g347(.A(G20), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n685), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n774), .C1(new_n611), .C2(new_n679), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n761), .A2(new_n762), .A3(new_n765), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n754), .A2(new_n755), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT98), .ZN(new_n780));
  INV_X1    g355(.A(G32), .ZN(new_n781));
  AOI21_X1  g356(.A(KEYINPUT96), .B1(new_n706), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n486), .A2(G141), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n483), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n479), .A2(G105), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n783), .A2(new_n784), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n706), .ZN(new_n789));
  MUX2_X1   g364(.A(new_n782), .B(KEYINPUT96), .S(new_n789), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n706), .A2(G26), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n486), .A2(KEYINPUT92), .A3(G140), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n795));
  INV_X1    g370(.A(G140), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n485), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n794), .A2(new_n797), .B1(G128), .B2(new_n483), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n793), .B1(new_n802), .B2(new_n706), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n793), .B(new_n803), .S(KEYINPUT28), .Z(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT24), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n706), .B1(new_n807), .B2(G34), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT94), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(G34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(KEYINPUT94), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G160), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n706), .ZN(new_n814));
  INV_X1    g389(.A(G2084), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT31), .B(G11), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  INV_X1    g393(.A(new_n628), .ZN(new_n819));
  INV_X1    g394(.A(G28), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT30), .ZN(new_n821));
  AOI21_X1  g396(.A(G29), .B1(new_n820), .B2(KEYINPUT30), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n819), .A2(G29), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n679), .A2(G21), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G168), .B2(new_n679), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1966), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n824), .B(new_n827), .C1(new_n746), .C2(new_n747), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n780), .A2(new_n792), .A3(new_n806), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n778), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n731), .A2(new_n732), .A3(new_n737), .A4(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n567), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G651), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(KEYINPUT99), .A3(G651), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n838), .A2(new_n839), .B1(G55), .B2(new_n527), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n534), .A2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n606), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT39), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n554), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT100), .B1(new_n550), .B2(new_n553), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n842), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n840), .A2(new_n849), .A3(new_n554), .A4(new_n841), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n848), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n844), .B1(new_n855), .B2(G860), .ZN(G145));
  XNOR2_X1  g431(.A(new_n713), .B(new_n621), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n483), .A2(G130), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n486), .A2(G142), .ZN(new_n859));
  NOR2_X1   g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(new_n469), .B2(G118), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n744), .A2(new_n801), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n503), .A2(new_n505), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(KEYINPUT4), .B2(new_n496), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n866), .A2(KEYINPUT102), .A3(new_n495), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n509), .B2(new_n510), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AND4_X1   g445(.A1(new_n739), .A2(new_n801), .A3(new_n741), .A4(new_n743), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n864), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n788), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n870), .B1(new_n864), .B2(new_n871), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n863), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n788), .ZN(new_n880));
  INV_X1    g455(.A(new_n863), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n875), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n628), .B(new_n813), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n490), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n881), .B1(new_n880), .B2(new_n875), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n882), .B1(new_n878), .B2(KEYINPUT103), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n886), .B(new_n887), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g469(.A1(G303), .A2(new_n681), .ZN(new_n895));
  NOR2_X1   g470(.A1(G166), .A2(G288), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G305), .ZN(new_n898));
  XOR2_X1   g473(.A(G290), .B(KEYINPUT105), .Z(new_n899));
  OAI21_X1  g474(.A(new_n694), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT107), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(KEYINPUT107), .B2(new_n906), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n854), .B(new_n616), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n606), .A2(G299), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n605), .A2(new_n611), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n606), .A2(KEYINPUT104), .A3(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n912), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n909), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n915), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n909), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n908), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n908), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n842), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n926), .ZN(G295));
  OAI21_X1  g502(.A(new_n925), .B1(G868), .B2(new_n926), .ZN(G331));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(G168), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(G286), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n853), .A3(new_n852), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n853), .B2(new_n852), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n918), .B1(new_n913), .B2(new_n914), .ZN(new_n936));
  INV_X1    g511(.A(new_n919), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n854), .A2(new_n930), .A3(new_n931), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n921), .A2(new_n939), .A3(new_n933), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n903), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n929), .B1(new_n941), .B2(G37), .ZN(new_n942));
  INV_X1    g517(.A(new_n903), .ZN(new_n943));
  INV_X1    g518(.A(new_n940), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n916), .A2(new_n919), .B1(new_n939), .B2(new_n933), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(KEYINPUT108), .A3(new_n887), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n938), .A2(new_n903), .A3(new_n940), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n942), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n918), .B1(new_n939), .B2(new_n933), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n917), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(new_n943), .C1(new_n921), .C2(new_n951), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n887), .A3(new_n949), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n955), .A3(KEYINPUT44), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n942), .A2(new_n947), .A3(new_n949), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n958), .A2(new_n959), .B1(KEYINPUT44), .B2(new_n962), .ZN(G397));
  XNOR2_X1  g538(.A(new_n801), .B(new_n805), .ZN(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n788), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n713), .A2(new_n716), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n717), .B2(new_n714), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n870), .B2(G1384), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT110), .B(G40), .ZN(new_n973));
  AND4_X1   g548(.A1(new_n477), .A2(new_n470), .A3(new_n480), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n970), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  NOR2_X1   g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n976), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n964), .A2(new_n968), .A3(new_n966), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n802), .A2(new_n805), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n873), .B2(new_n964), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n976), .A2(new_n965), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT46), .Z(new_n990));
  OR3_X1    g565(.A1(new_n988), .A2(KEYINPUT47), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT47), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n982), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT73), .B1(new_n866), .B2(new_n495), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n509), .A2(new_n508), .A3(new_n510), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n971), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT45), .B(new_n998), .C1(new_n867), .C2(new_n869), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n974), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1971), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n997), .A2(new_n1006), .A3(new_n998), .A4(new_n999), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n866), .A2(new_n495), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT50), .B1(new_n1008), .B2(G1384), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1007), .A2(new_n974), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n755), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n996), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G166), .A2(new_n996), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT55), .Z(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n995), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1004), .A2(new_n1003), .B1(new_n1010), .B2(new_n755), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT115), .B(new_n1014), .C1(new_n1017), .C2(new_n996), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1006), .B(new_n998), .C1(new_n866), .C2(new_n495), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n974), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(KEYINPUT50), .B2(new_n1000), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n755), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1005), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(G8), .A3(new_n1015), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT112), .B1(new_n694), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n1029));
  NOR4_X1   g604(.A1(new_n690), .A2(new_n693), .A3(new_n1029), .A4(G1981), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT49), .B(new_n1026), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT113), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1026), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n509), .B2(new_n510), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n996), .B1(new_n1036), .B2(new_n974), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1029), .B1(G305), .B2(G1981), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n694), .A2(KEYINPUT112), .A3(new_n1027), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT49), .A4(new_n1026), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n681), .A2(G1976), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1037), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G288), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(KEYINPUT111), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1037), .A2(new_n1046), .A3(new_n1048), .A4(new_n1044), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1046), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1043), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT116), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1043), .A2(new_n1049), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1021), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n815), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n971), .B1(new_n1008), .B2(G1384), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n974), .B(new_n1063), .C1(new_n1000), .C2(new_n971), .ZN(new_n1064));
  INV_X1    g639(.A(G1966), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1022), .A2(new_n1067), .A3(new_n815), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G8), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(G286), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1019), .A2(new_n1025), .A3(new_n1058), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1024), .A2(G8), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1075), .B2(new_n1014), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1054), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1071), .A2(new_n1076), .A3(new_n1025), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G168), .A2(new_n996), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n1081), .B2(KEYINPUT124), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1069), .A2(G8), .A3(G286), .ZN(new_n1085));
  OAI211_X1 g660(.A(G8), .B(new_n1082), .C1(new_n1069), .C2(G286), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT62), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n996), .B(new_n1014), .C1(new_n1005), .C2(new_n1023), .ZN(new_n1089));
  AOI221_X4 g664(.A(new_n1089), .B1(new_n1055), .B2(new_n1057), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1003), .B2(G2078), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1006), .B1(new_n512), .B2(new_n998), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n769), .B1(new_n1093), .B2(new_n1021), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1064), .A2(new_n1091), .A3(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1084), .A2(new_n1098), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1088), .A2(new_n1090), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1025), .A2(new_n1054), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1036), .A2(new_n974), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1043), .A2(new_n1047), .A3(new_n681), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n996), .B(new_n1103), .C1(new_n1104), .C2(new_n1040), .ZN(new_n1105));
  OR3_X1    g680(.A1(new_n1101), .A2(new_n1105), .A3(KEYINPUT114), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT114), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1079), .A2(new_n1100), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1007), .A2(new_n974), .A3(new_n1009), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1001), .A2(new_n974), .A3(new_n1002), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(KEYINPUT118), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n611), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1118), .A3(KEYINPUT57), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n573), .B2(new_n575), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n610), .A2(new_n572), .A3(KEYINPUT118), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1115), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1102), .A2(G2067), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1022), .B2(G1348), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n605), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1132), .A2(new_n1136), .B1(new_n1138), .B2(new_n1135), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1001), .A2(new_n965), .A3(new_n1002), .A4(new_n974), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1102), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n554), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n554), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1143), .A2(new_n1149), .A3(new_n554), .A4(new_n1144), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1139), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1129), .A2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g729(.A(KEYINPUT122), .B(new_n605), .C1(new_n1129), .C2(new_n1153), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1348), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1153), .B1(new_n1157), .B2(new_n1127), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1158), .B2(new_n606), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1154), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n759), .B1(new_n1093), .B2(new_n1021), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT60), .B1(new_n1161), .B2(new_n1128), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT122), .B1(new_n1162), .B2(new_n605), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1154), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(new_n1156), .A3(new_n606), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(KEYINPUT123), .B(new_n1134), .C1(new_n1152), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1155), .A2(new_n1159), .A3(new_n1154), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1164), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1151), .B(new_n1139), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1172), .B2(new_n1133), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1002), .A2(G160), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1091), .A2(G2078), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(G40), .A3(new_n972), .A4(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1095), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1097), .B1(G301), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1087), .B1(new_n1179), .B2(KEYINPUT54), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1092), .A2(new_n1177), .A3(new_n1094), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(G171), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1182), .A2(KEYINPUT125), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT54), .B1(new_n1182), .B2(KEYINPUT125), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1095), .A2(G301), .A3(new_n1096), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1090), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1180), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1109), .B1(new_n1174), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n970), .B1(G1986), .B2(G290), .ZN(new_n1190));
  INV_X1    g765(.A(new_n979), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n983), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n994), .B1(new_n1189), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g768(.A(G227), .B1(G14), .B2(new_n644), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n893), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G229), .A2(new_n465), .ZN(new_n1197));
  INV_X1    g771(.A(new_n1197), .ZN(new_n1198));
  NOR3_X1   g772(.A1(new_n1196), .A2(new_n962), .A3(new_n1198), .ZN(G308));
  NOR2_X1   g773(.A1(new_n962), .A2(new_n1198), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1200), .A2(new_n893), .A3(new_n1195), .ZN(G225));
endmodule


