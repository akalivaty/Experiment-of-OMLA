//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G190gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n204), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n215), .A2(new_n216), .A3(new_n211), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n215), .B2(new_n211), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(KEYINPUT26), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n221), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n231), .A2(new_n233), .A3(new_n235), .A4(new_n224), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n230), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n231), .A2(new_n235), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n221), .A2(new_n237), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n233), .A2(new_n224), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(KEYINPUT25), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n219), .A2(new_n229), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n202), .B1(new_n244), .B2(KEYINPUT29), .ZN(new_n245));
  INV_X1    g044(.A(new_n229), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n215), .A2(new_n211), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n216), .A3(new_n211), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n250), .B2(new_n213), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n239), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(G226gat), .B(G233gat), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n261), .B(new_n255), .C1(new_n258), .C2(new_n259), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n245), .A2(new_n254), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT70), .B(KEYINPUT29), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n202), .B1(new_n244), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT71), .B(new_n202), .C1(new_n244), .C2(new_n268), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n254), .ZN(new_n273));
  INV_X1    g072(.A(new_n265), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT72), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n254), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n267), .B1(new_n251), .B2(new_n253), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n282), .B2(new_n202), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n274), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n266), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n278), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n285), .A3(new_n279), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT30), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n292), .A3(new_n279), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(G134gat), .ZN(new_n299));
  INV_X1    g098(.A(G134gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G127gat), .ZN(new_n301));
  OAI22_X1  g100(.A1(new_n297), .A2(KEYINPUT1), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G134gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n317), .A2(KEYINPUT74), .B1(KEYINPUT2), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G155gat), .B(G162gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT73), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(G162gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G155gat), .ZN(new_n326));
  OR2_X1    g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n326), .A2(KEYINPUT2), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n314), .A2(KEYINPUT75), .ZN(new_n329));
  MUX2_X1   g128(.A(KEYINPUT75), .B(new_n329), .S(new_n316), .Z(new_n330));
  AOI22_X1  g129(.A1(new_n322), .A2(new_n324), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n312), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n322), .A2(new_n324), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n328), .A2(new_n330), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n296), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n335), .A3(new_n311), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n339), .A2(KEYINPUT78), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT78), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n334), .A2(new_n335), .A3(new_n345), .A4(new_n311), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n296), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n334), .A2(new_n335), .A3(new_n311), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n311), .B1(new_n334), .B2(new_n335), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(KEYINPUT80), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT5), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n334), .A2(new_n335), .A3(new_n311), .A4(new_n340), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n331), .A2(KEYINPUT83), .A3(new_n311), .A4(new_n340), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n331), .A2(new_n332), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n312), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n368));
  OAI22_X1  g167(.A1(new_n349), .A2(new_n357), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G1gat), .B(G29gat), .Z(new_n370));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT82), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n372), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(new_n350), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n351), .A2(new_n352), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n296), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT39), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n296), .B1(new_n363), .B2(new_n366), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT39), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n383), .A2(KEYINPUT40), .A3(new_n375), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT40), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n375), .B1(new_n384), .B2(new_n381), .ZN(new_n389));
  AOI211_X1 g188(.A(KEYINPUT39), .B(new_n296), .C1(new_n363), .C2(new_n366), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n377), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n295), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n394), .B(KEYINPUT85), .Z(new_n395));
  AOI21_X1  g194(.A(new_n265), .B1(new_n365), .B2(new_n267), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n267), .B1(new_n262), .B2(new_n264), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n331), .B1(new_n397), .B2(new_n332), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n262), .B2(new_n264), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n401), .A2(KEYINPUT86), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT3), .B1(new_n401), .B2(KEYINPUT86), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n331), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n268), .B1(new_n331), .B2(new_n332), .ZN(new_n405));
  OAI211_X1 g204(.A(G228gat), .B(G233gat), .C1(new_n405), .C2(new_n265), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n399), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G22gat), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n399), .B(new_n409), .C1(new_n404), .C2(new_n406), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT84), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n411), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT38), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n286), .A2(KEYINPUT37), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n279), .B1(new_n286), .B2(KEYINPUT37), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(KEYINPUT87), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n278), .B1(new_n275), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n417), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  OAI221_X1 g225(.A(new_n375), .B1(new_n367), .B2(new_n368), .C1(new_n349), .C2(new_n357), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n377), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n369), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n278), .A2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n273), .A2(new_n265), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n245), .A2(new_n254), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n421), .B1(new_n432), .B2(new_n274), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(KEYINPUT37), .B2(new_n286), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n428), .A2(new_n429), .A3(new_n290), .A4(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n393), .B(new_n416), .C1(new_n425), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n411), .B(new_n414), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n428), .A2(new_n429), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n440), .B2(new_n295), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442));
  AOI221_X4 g241(.A(new_n311), .B1(new_n239), .B2(new_n243), .C1(new_n219), .C2(new_n229), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n219), .A2(new_n229), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n312), .B1(new_n444), .B2(new_n252), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G227gat), .ZN(new_n447));
  INV_X1    g246(.A(G233gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT67), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT67), .ZN(new_n451));
  INV_X1    g250(.A(new_n449), .ZN(new_n452));
  NOR4_X1   g251(.A1(new_n443), .A2(new_n445), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n442), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT32), .B1(new_n450), .B2(new_n453), .ZN(new_n455));
  XOR2_X1   g254(.A(G15gat), .B(G43gat), .Z(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n452), .B1(new_n443), .B2(new_n445), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n458), .ZN(new_n464));
  OAI221_X1 g263(.A(KEYINPUT32), .B1(new_n442), .B2(new_n464), .C1(new_n450), .C2(new_n453), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n459), .A2(KEYINPUT68), .A3(new_n463), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n463), .B1(new_n459), .B2(new_n465), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT36), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n474), .B(new_n471), .C1(new_n468), .C2(new_n469), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n437), .B(new_n441), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n416), .A3(new_n472), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n280), .A2(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n479));
  NAND2_X1  g278(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n439), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n477), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n481), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n471), .B1(new_n468), .B2(new_n469), .ZN(new_n484));
  INV_X1    g283(.A(new_n477), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n483), .A2(new_n416), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n476), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT16), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(G1gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  MUX2_X1   g289(.A(G1gat), .B(new_n489), .S(new_n490), .Z(new_n491));
  XOR2_X1   g290(.A(new_n491), .B(G8gat), .Z(new_n492));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  INV_X1    g293(.A(G36gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n496), .A2(new_n497), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n499), .B2(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n500), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n499), .A2(new_n504), .A3(KEYINPUT15), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(KEYINPUT91), .A3(new_n498), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n498), .A3(new_n507), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n503), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n492), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(KEYINPUT17), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n503), .A2(new_n511), .A3(new_n515), .A4(new_n508), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n492), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT18), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT92), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n519), .A2(new_n523), .A3(KEYINPUT18), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT18), .B1(new_n519), .B2(new_n520), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n492), .B(new_n512), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n520), .B(KEYINPUT13), .Z(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT11), .ZN(new_n531));
  INV_X1    g330(.A(G169gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G197gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT12), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n526), .B2(KEYINPUT93), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n525), .A2(new_n529), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n525), .B2(new_n529), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542));
  MUX2_X1   g341(.A(KEYINPUT7), .B(new_n541), .S(new_n542), .Z(new_n543));
  INV_X1    g342(.A(KEYINPUT8), .ZN(new_n544));
  INV_X1    g343(.A(G99gat), .ZN(new_n545));
  INV_X1    g344(.A(G106gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT97), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(G99gat), .A3(G106gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n543), .A2(new_n550), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n517), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n512), .A2(new_n557), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n559), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n557), .B1(new_n514), .B2(new_n516), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n568), .B2(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n567), .B(new_n569), .C1(KEYINPUT41), .C2(new_n561), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G134gat), .B(G162gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  INV_X1    g376(.A(G57gat), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT94), .B1(new_n578), .B2(G64gat), .ZN(new_n579));
  INV_X1    g378(.A(G64gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G57gat), .ZN(new_n581));
  MUX2_X1   g380(.A(KEYINPUT94), .B(new_n579), .S(new_n581), .Z(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(KEYINPUT9), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n581), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n580), .A2(G57gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT9), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n585), .A2(new_n586), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n518), .B1(new_n577), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT96), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G231gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n448), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n594), .B2(new_n577), .ZN(new_n602));
  AOI211_X1 g401(.A(KEYINPUT21), .B(new_n600), .C1(new_n588), .C2(new_n593), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n582), .A2(new_n587), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n591), .B2(new_n592), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n600), .B1(new_n606), .B2(KEYINPUT21), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n594), .A2(new_n577), .A3(new_n601), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n597), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT95), .Z(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n604), .B2(new_n609), .ZN(new_n614));
  XOR2_X1   g413(.A(G183gat), .B(G211gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n604), .A2(new_n609), .ZN(new_n618));
  INV_X1    g417(.A(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n620), .B2(new_n612), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n596), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n596), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n612), .A3(new_n615), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n616), .B1(new_n613), .B2(new_n614), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n575), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n572), .A2(new_n573), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n576), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n553), .B1(new_n555), .B2(KEYINPUT98), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n551), .A2(new_n635), .A3(new_n552), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n594), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n554), .A2(new_n556), .B1(new_n588), .B2(new_n593), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n557), .A2(new_n606), .A3(KEYINPUT10), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n632), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n634), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n606), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n557), .A2(new_n594), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT10), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n631), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n645), .A3(new_n632), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n642), .A2(new_n650), .A3(new_n651), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n651), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT100), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n540), .A2(new_n630), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n487), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n439), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n479), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(G8gat), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n671), .B(new_n673), .C1(KEYINPUT42), .C2(new_n672), .ZN(G1325gat));
  NOR2_X1   g473(.A1(new_n473), .A2(new_n475), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n665), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n484), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n665), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n416), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n576), .A2(new_n629), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n487), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n525), .A2(new_n529), .ZN(new_n686));
  INV_X1    g485(.A(new_n537), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n525), .A2(new_n529), .A3(new_n537), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n663), .ZN(new_n691));
  INV_X1    g490(.A(new_n627), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n494), .A3(new_n440), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT102), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n487), .A2(KEYINPUT44), .A3(new_n684), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n487), .B2(new_n684), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n701), .A3(new_n693), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n699), .B1(new_n703), .B2(new_n439), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(KEYINPUT103), .A3(new_n440), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(G29gat), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n696), .A2(new_n697), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n698), .A2(new_n706), .A3(new_n707), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n694), .A2(new_n495), .A3(new_n295), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n703), .B2(new_n479), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n702), .A2(new_n675), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n702), .A2(KEYINPUT104), .A3(new_n675), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n678), .A2(G43gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n694), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT47), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n714), .A2(G43gat), .B1(new_n694), .B2(new_n719), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n718), .A2(new_n721), .B1(new_n722), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g522(.A1(new_n702), .A2(G50gat), .A3(new_n438), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n685), .A2(new_n416), .A3(new_n693), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(G50gat), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n690), .A2(new_n630), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n691), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n487), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n439), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT105), .B(G57gat), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1332gat));
  INV_X1    g533(.A(new_n731), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n735), .B(new_n295), .C1(new_n736), .C2(new_n580), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT106), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n580), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  NOR2_X1   g539(.A1(new_n731), .A2(new_n678), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT107), .B1(new_n731), .B2(new_n678), .ZN(new_n744));
  AOI21_X1  g543(.A(G71gat), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n583), .B1(new_n735), .B2(new_n675), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT109), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n744), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n731), .A2(KEYINPUT107), .A3(new_n678), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n583), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  INV_X1    g550(.A(new_n746), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n747), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n747), .B2(new_n753), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1334gat));
  NOR2_X1   g556(.A1(new_n731), .A2(new_n416), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n584), .ZN(G1335gat));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n690), .A2(new_n627), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n663), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n700), .A2(new_n701), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n760), .B1(new_n764), .B2(new_n439), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(KEYINPUT110), .A3(new_n440), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(G85gat), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n476), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n482), .A2(new_n486), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n684), .B(new_n761), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n487), .A2(KEYINPUT51), .A3(new_n684), .A4(new_n761), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n691), .A2(G85gat), .A3(new_n439), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(G92gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n763), .B2(new_n295), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n770), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n770), .B2(KEYINPUT111), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n691), .A2(G92gat), .A3(new_n479), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n786));
  AND2_X1   g585(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n775), .A2(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n779), .B2(new_n788), .ZN(G1337gat));
  OAI21_X1  g588(.A(G99gat), .B1(new_n764), .B2(new_n676), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n484), .A2(new_n545), .A3(new_n663), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n775), .B2(new_n791), .ZN(G1338gat));
  AOI21_X1  g591(.A(new_n546), .B1(new_n763), .B2(new_n438), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n691), .A2(G106gat), .A3(new_n416), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n781), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n685), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n487), .A2(KEYINPUT44), .A3(new_n684), .ZN(new_n800));
  INV_X1    g599(.A(new_n762), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n799), .A2(new_n438), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT53), .B1(new_n802), .B2(G106gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n774), .B2(new_n794), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT113), .B(new_n795), .C1(new_n772), .C2(new_n773), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n797), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n729), .A2(new_n663), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n519), .A2(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n814));
  INV_X1    g613(.A(new_n535), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n536), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n525), .A2(new_n529), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n663), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n655), .B1(new_n641), .B2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n646), .A2(new_n647), .A3(new_n631), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n642), .A2(new_n650), .A3(KEYINPUT54), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT55), .B(new_n821), .C1(new_n823), .C2(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n656), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n819), .B1(new_n540), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n684), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n829), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n684), .A3(new_n816), .A4(new_n818), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n813), .B1(new_n835), .B2(new_n692), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n439), .A2(new_n295), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n416), .A3(new_n484), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n305), .B1(new_n840), .B2(new_n540), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n836), .B2(new_n438), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n627), .B1(new_n832), .B2(new_n834), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT116), .B(new_n416), .C1(new_n844), .C2(new_n813), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n484), .A3(new_n837), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n690), .A2(G113gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n841), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT117), .ZN(G1340gat));
  NOR3_X1   g649(.A1(new_n847), .A2(new_n303), .A3(new_n691), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n840), .A2(new_n691), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n303), .B2(new_n852), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n847), .B2(new_n692), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n627), .A2(new_n298), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n840), .B2(new_n855), .ZN(G1342gat));
  NOR2_X1   g655(.A1(new_n836), .A2(new_n439), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n684), .A2(new_n479), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT118), .Z(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(G134gat), .A3(new_n478), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT56), .Z(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n847), .B2(new_n831), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n676), .A2(new_n837), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n836), .B2(new_n416), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n438), .C1(new_n844), .C2(new_n813), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n313), .B1(new_n869), .B2(new_n690), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n675), .A2(new_n416), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n839), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(G141gat), .A3(new_n540), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n870), .A2(KEYINPUT58), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT58), .B1(new_n870), .B2(new_n873), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1344gat));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n728), .B2(new_n691), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n690), .A2(new_n630), .A3(new_n663), .A4(KEYINPUT121), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n438), .B1(new_n844), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n868), .A2(new_n878), .B1(new_n883), .B2(new_n866), .ZN(new_n884));
  INV_X1    g683(.A(new_n836), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n438), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n865), .B(KEYINPUT119), .Z(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n663), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n877), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT59), .B(new_n315), .C1(new_n869), .C2(new_n663), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n857), .A2(new_n871), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n663), .A2(new_n315), .A3(new_n479), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(new_n893), .ZN(G1345gat));
  NOR2_X1   g693(.A1(new_n872), .A2(new_n692), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n896));
  AOI21_X1  g695(.A(G155gat), .B1(new_n895), .B2(KEYINPUT122), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n627), .A2(G155gat), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(new_n869), .B2(new_n898), .ZN(G1346gat));
  OR3_X1    g698(.A1(new_n892), .A2(new_n325), .A3(new_n859), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n869), .A2(new_n684), .ZN(new_n901));
  INV_X1    g700(.A(new_n325), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G1347gat));
  NOR4_X1   g702(.A1(new_n836), .A2(new_n440), .A3(new_n479), .A4(new_n478), .ZN(new_n904));
  AOI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n690), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n440), .A2(new_n479), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n678), .B(new_n908), .C1(new_n843), .C2(new_n845), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n540), .A2(new_n532), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n846), .A2(new_n484), .A3(new_n907), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n912), .B2(new_n691), .ZN(new_n913));
  INV_X1    g712(.A(G176gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n904), .A2(new_n914), .A3(new_n663), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1349gat));
  AOI21_X1  g715(.A(new_n203), .B1(new_n909), .B2(new_n627), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n904), .A2(new_n208), .A3(new_n210), .A4(new_n627), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT60), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G183gat), .B1(new_n912), .B2(new_n692), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n214), .A3(new_n684), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n846), .A2(new_n484), .A3(new_n684), .A4(new_n907), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(G190gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n926), .B2(G190gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n836), .A2(new_n440), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n871), .A2(new_n295), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n690), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n907), .A2(new_n676), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT125), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n884), .B2(new_n886), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n540), .A2(new_n534), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(new_n939), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n887), .A2(new_n663), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n946), .A3(new_n663), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(G204gat), .A3(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n935), .A2(G204gat), .A3(new_n691), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1353gat));
  OR3_X1    g750(.A1(new_n935), .A2(G211gat), .A3(new_n692), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n907), .A2(new_n676), .A3(new_n627), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n887), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n684), .B1(new_n940), .B2(new_n959), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT127), .B(new_n939), .C1(new_n884), .C2(new_n886), .ZN(new_n961));
  OAI21_X1  g760(.A(G218gat), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n935), .A2(G218gat), .A3(new_n831), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


