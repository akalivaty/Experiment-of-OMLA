//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n203), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n221));
  AND3_X1   g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n218), .A2(new_n222), .B1(G1), .B2(G20), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n216), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(new_n224), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n238), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  AND3_X1   g0046(.A1(new_n246), .A2(KEYINPUT68), .A3(new_n213), .ZN(new_n247));
  AOI21_X1  g0047(.A(KEYINPUT68), .B1(new_n246), .B2(new_n213), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G50), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n214), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n214), .A2(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G58), .A2(G68), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n214), .B1(new_n262), .B2(new_n239), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n249), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n252), .A2(new_n239), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n255), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n213), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n270), .A2(KEYINPUT66), .A3(G222), .A4(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT66), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n278), .B2(G77), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n272), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(new_n278), .B2(new_n271), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n270), .A2(KEYINPUT67), .A3(G1698), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n269), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n291), .A3(G274), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(G226), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n286), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G169), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n267), .B(new_n300), .C1(new_n301), .C2(new_n299), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(KEYINPUT69), .A3(G190), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n298), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n255), .A2(new_n311), .A3(new_n264), .A4(new_n265), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n310), .A2(new_n312), .B1(new_n298), .B2(G200), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n308), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n308), .B2(new_n313), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n303), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n251), .A2(KEYINPUT70), .A3(G68), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT12), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT70), .B1(new_n251), .B2(G68), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G20), .A2(G33), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n257), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n249), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n321), .B(new_n322), .C1(new_n323), .C2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n253), .A2(G68), .A3(new_n254), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n323), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n275), .A2(new_n277), .A3(G232), .A4(G1698), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(new_n271), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n269), .ZN(new_n340));
  INV_X1    g0140(.A(G274), .ZN(new_n341));
  AND2_X1   g0141(.A1(G1), .A2(G13), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n290), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n296), .A2(G238), .B1(new_n289), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n340), .B2(new_n344), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n335), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n344), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(G179), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n335), .B1(new_n354), .B2(G169), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n334), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(G200), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n333), .C1(new_n306), .C2(new_n354), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n256), .B1(new_n250), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n253), .A2(new_n360), .B1(new_n252), .B2(new_n256), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n246), .A2(new_n213), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n246), .A2(KEYINPUT68), .A3(new_n213), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n270), .B2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n214), .B1(new_n203), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G159), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n260), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n373), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n262), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n324), .A2(G159), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(KEYINPUT71), .A3(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n371), .A2(G68), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n367), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n202), .B1(new_n369), .B2(new_n370), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n379), .A2(new_n380), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n362), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n292), .B1(new_n228), .B2(new_n295), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n275), .A2(new_n277), .A3(G223), .A4(new_n271), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n269), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G169), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n269), .B2(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G179), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n388), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n371), .A2(G68), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n377), .A2(new_n381), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n249), .A3(new_n387), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n361), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n397), .A2(new_n399), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n390), .A2(new_n395), .A3(new_n306), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n398), .B2(G200), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n411), .A3(new_n361), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n405), .A2(new_n411), .A3(KEYINPUT17), .A4(new_n361), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n401), .A2(new_n409), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n293), .B1(G244), .B2(new_n296), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n270), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n283), .A2(new_n284), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(G238), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n418), .B1(new_n423), .B2(new_n291), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n306), .ZN(new_n425));
  INV_X1    g0225(.A(new_n256), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n324), .B1(G20), .B2(G77), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT15), .B(G87), .Z(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n257), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n249), .B1(new_n326), .B2(new_n252), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n253), .A2(G77), .A3(new_n254), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n424), .A2(G200), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G169), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n301), .B(new_n418), .C1(new_n423), .C2(new_n291), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n359), .A2(new_n417), .A3(new_n436), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n316), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n288), .A2(G1), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n291), .A2(G274), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n250), .A2(G45), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(G250), .C1(new_n268), .C2(new_n213), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n275), .A2(new_n277), .A3(G238), .A4(new_n271), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n451), .B2(new_n269), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G190), .ZN(new_n453));
  INV_X1    g0253(.A(G200), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n452), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n428), .A2(new_n251), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT19), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n214), .B1(new_n338), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G87), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n420), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n275), .A2(new_n277), .A3(new_n214), .A4(G68), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n457), .B1(new_n257), .B2(new_n460), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n456), .B1(new_n465), .B2(new_n249), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n250), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n367), .A2(G87), .A3(new_n251), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n367), .A2(new_n251), .A3(new_n428), .A4(new_n467), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n451), .A2(new_n269), .ZN(new_n472));
  INV_X1    g0272(.A(new_n447), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n301), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n452), .A2(G169), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n455), .A2(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n275), .A2(new_n277), .A3(new_n214), .A4(G87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT22), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n270), .A2(new_n480), .A3(new_n214), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n420), .A3(G20), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT80), .A2(KEYINPUT24), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n482), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n491), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n493), .B(new_n488), .C1(new_n479), .C2(new_n481), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n249), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND4_X1   g0295(.A1(G107), .A2(new_n367), .A3(new_n251), .A4(new_n467), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n252), .A2(new_n420), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT74), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT73), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n287), .A3(KEYINPUT5), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(KEYINPUT73), .B2(G41), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n505), .A3(new_n443), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n291), .A2(G274), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n287), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n445), .B1(new_n509), .B2(new_n504), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(KEYINPUT74), .A3(new_n343), .A4(new_n503), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n269), .B1(new_n510), .B2(new_n503), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G264), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(new_n271), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n269), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n512), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G179), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n437), .B2(new_n520), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n477), .B1(new_n500), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n420), .B1(new_n369), .B2(new_n370), .ZN(new_n524));
  AND4_X1   g0324(.A1(KEYINPUT72), .A2(new_n214), .A3(new_n259), .A4(G77), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT72), .B1(new_n324), .B2(G77), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT6), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n214), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n249), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n253), .A2(G97), .A3(new_n467), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n252), .A2(new_n460), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT75), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(new_n539), .A3(new_n535), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n508), .A2(new_n511), .B1(new_n513), .B2(G257), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(new_n271), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n543), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n269), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n437), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n542), .A2(G179), .A3(new_n549), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n547), .ZN(new_n555));
  INV_X1    g0355(.A(new_n548), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n291), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n513), .A2(G257), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n512), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n557), .A2(new_n559), .A3(new_n306), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n454), .B1(new_n542), .B2(new_n549), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n560), .A2(new_n537), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n520), .A2(G190), .ZN(new_n564));
  AOI22_X1  g0364(.A1(G264), .A2(new_n513), .B1(new_n518), .B2(new_n269), .ZN(new_n565));
  AOI21_X1  g0365(.A(G200), .B1(new_n565), .B2(new_n512), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n495), .B(new_n499), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n523), .A2(new_n554), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n513), .A2(G270), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n276), .A2(G33), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n571));
  OAI21_X1  g0371(.A(G303), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n275), .A2(new_n277), .A3(G264), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(new_n271), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n269), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n512), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n543), .B(new_n214), .C1(G33), .C2(new_n460), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G20), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n363), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n363), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n367), .A2(G116), .A3(new_n251), .A4(new_n467), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n252), .A2(new_n579), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n577), .A2(new_n588), .A3(G169), .ZN(new_n589));
  XNOR2_X1  g0389(.A(KEYINPUT77), .B(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(KEYINPUT78), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT79), .ZN(new_n596));
  AOI22_X1  g0396(.A1(G270), .A2(new_n513), .B1(new_n575), .B2(new_n269), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n454), .B1(new_n597), .B2(new_n512), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n598), .B2(new_n588), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n577), .A2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(new_n588), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(KEYINPUT79), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n599), .B(new_n602), .C1(new_n306), .C2(new_n577), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n512), .A2(new_n569), .A3(new_n576), .A4(G179), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n577), .A2(new_n588), .A3(KEYINPUT21), .A4(G169), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT76), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n437), .B1(new_n597), .B2(new_n512), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT76), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT21), .A4(new_n588), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n595), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n568), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n442), .A2(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n414), .A2(new_n415), .ZN(new_n615));
  INV_X1    g0415(.A(new_n440), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n358), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n615), .B1(new_n617), .B2(new_n356), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n401), .A2(new_n409), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n314), .A2(new_n315), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n303), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT83), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT83), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n303), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n469), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n453), .C1(new_n454), .C2(new_n452), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n301), .A2(new_n452), .B1(new_n466), .B2(new_n470), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n472), .A2(new_n473), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT81), .B1(new_n630), .B2(new_n437), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT81), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n452), .A2(new_n632), .A3(G169), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n629), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n567), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n538), .A2(new_n540), .B1(new_n551), .B2(new_n552), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(new_n562), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n595), .A2(new_n611), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT82), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT82), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n595), .A2(new_n611), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n521), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n520), .A2(new_n437), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n500), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n638), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n634), .A2(new_n628), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(new_n552), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n537), .B1(new_n651), .B2(new_n550), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n634), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n306), .B(new_n447), .C1(new_n269), .C2(new_n451), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n454), .B1(new_n472), .B2(new_n473), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n630), .A2(new_n437), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n658), .A2(new_n627), .B1(new_n629), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n650), .B1(new_n636), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n442), .B1(new_n647), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n626), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(new_n646), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n250), .A2(new_n214), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n567), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n500), .B2(new_n672), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n666), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT84), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n601), .A2(new_n673), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n640), .A2(new_n642), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n612), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n639), .A2(new_n673), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n678), .A2(new_n687), .B1(new_n666), .B2(new_n673), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n461), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n211), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n648), .B2(new_n652), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n541), .A2(new_n650), .A3(new_n660), .A4(new_n553), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n634), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT86), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT86), .A4(new_n634), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n595), .A2(new_n611), .A3(new_n646), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n637), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n697), .B1(new_n706), .B2(new_n673), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n520), .B1(new_n557), .B2(new_n559), .ZN(new_n709));
  AOI21_X1  g0509(.A(G179), .B1(new_n472), .B2(new_n473), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n577), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT30), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n542), .A2(new_n565), .A3(new_n549), .A4(new_n452), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(KEYINPUT85), .B2(new_n604), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT85), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n597), .A2(new_n715), .A3(G179), .A4(new_n512), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n577), .A2(new_n710), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n549), .A2(new_n542), .B1(new_n565), .B2(new_n512), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n604), .A2(KEYINPUT85), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n557), .A2(new_n559), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n565), .A2(new_n452), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n716), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n717), .A2(new_n726), .A3(new_n672), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n613), .B2(new_n673), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n708), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n595), .A2(new_n611), .A3(new_n641), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n641), .B1(new_n595), .B2(new_n611), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n646), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n637), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n672), .B1(new_n736), .B2(new_n662), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n707), .B(new_n732), .C1(new_n697), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT87), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n696), .B1(new_n739), .B2(G1), .ZN(G364));
  INV_X1    g0540(.A(new_n683), .ZN(new_n741));
  INV_X1    g0541(.A(G13), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n250), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n691), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n682), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n213), .B1(G20), .B2(new_n437), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT89), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT89), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT90), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n690), .A2(new_n270), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n244), .A2(new_n288), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n759), .B(new_n760), .C1(new_n288), .C2(new_n212), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n270), .A2(new_n207), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n207), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(KEYINPUT88), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(KEYINPUT88), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n757), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n746), .ZN(new_n768));
  NAND2_X1  g0568(.A1(G20), .A2(G179), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT91), .ZN(new_n770));
  AOI21_X1  g0570(.A(G200), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n306), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  INV_X1    g0575(.A(G326), .ZN(new_n776));
  NAND4_X1  g0576(.A1(G20), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT92), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n772), .A2(G190), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(G311), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n454), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G20), .A3(G190), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n278), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G20), .A3(new_n306), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n790), .B1(G329), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n214), .B1(new_n791), .B2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n769), .A2(new_n454), .A3(G190), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(G294), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(G20), .A3(new_n306), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n794), .B(new_n799), .C1(new_n800), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G107), .ZN(new_n807));
  OAI21_X1  g0607(.A(KEYINPUT32), .B1(new_n792), .B2(new_n375), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n788), .A2(new_n459), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n278), .B(new_n809), .C1(G68), .C2(new_n797), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n792), .A2(KEYINPUT32), .A3(new_n375), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G97), .B2(new_n796), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n782), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(G50), .B1(new_n784), .B2(G77), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n201), .B2(new_n774), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n786), .A2(new_n805), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT94), .ZN(new_n819));
  INV_X1    g0619(.A(new_n752), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n818), .B2(KEYINPUT94), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n767), .B(new_n768), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n755), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n682), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n748), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NOR2_X1   g0626(.A1(new_n752), .A2(new_n753), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n746), .B1(new_n828), .B2(G77), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n814), .A2(G137), .B1(new_n784), .B2(G159), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n773), .A2(G143), .B1(G150), .B2(new_n797), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n806), .A2(G68), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n270), .B1(new_n788), .B2(new_n239), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G132), .B2(new_n793), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n201), .C2(new_n795), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n804), .A2(new_n459), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n278), .B1(new_n792), .B2(new_n839), .C1(new_n788), .C2(new_n420), .ZN(new_n840));
  INV_X1    g0640(.A(new_n797), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n841), .A2(new_n800), .B1(new_n795), .B2(new_n460), .ZN(new_n842));
  OR3_X1    g0642(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G116), .A2(new_n784), .B1(new_n773), .B2(G294), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n789), .B2(new_n782), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n833), .A2(new_n837), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n829), .B1(new_n846), .B2(new_n752), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n433), .B(new_n672), .C1(new_n616), .C2(KEYINPUT95), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT95), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n433), .A2(new_n672), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n440), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n848), .A2(new_n851), .B1(new_n435), .B2(new_n434), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n847), .B1(new_n852), .B2(new_n754), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n737), .A2(new_n852), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n673), .B(new_n852), .C1(new_n647), .C2(new_n663), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n732), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT96), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n732), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n746), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n854), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n743), .A2(new_n250), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n619), .A2(new_n670), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT98), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n377), .A2(new_n381), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n385), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n402), .A2(KEYINPUT98), .A3(new_n403), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n384), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n362), .B1(new_n869), .B2(new_n383), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n412), .B1(new_n870), .B2(new_n400), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n670), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n406), .A2(new_n408), .ZN(new_n874));
  INV_X1    g0674(.A(new_n670), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n406), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n876), .A3(new_n412), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n416), .A2(KEYINPUT99), .A3(new_n872), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT99), .B1(new_n416), .B2(new_n872), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT38), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n874), .A2(new_n876), .A3(new_n412), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n877), .ZN(new_n888));
  INV_X1    g0688(.A(new_n876), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n416), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n883), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n886), .B1(KEYINPUT39), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n356), .A2(new_n672), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n864), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT101), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n416), .A2(new_n872), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT99), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n416), .A2(KEYINPUT99), .A3(new_n872), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n901), .B2(new_n879), .ZN(new_n902));
  INV_X1    g0702(.A(new_n885), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n896), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n885), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT97), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n353), .A2(new_n355), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n358), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n333), .A2(new_n673), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n910), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n356), .A2(new_n358), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AND4_X1   g0714(.A1(new_n907), .A2(new_n356), .A3(new_n358), .A4(new_n912), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n440), .A2(new_n672), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n856), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n895), .B1(new_n906), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n707), .B1(new_n737), .B2(new_n697), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n923), .A2(new_n442), .B1(new_n625), .B2(new_n623), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n921), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n727), .A2(KEYINPUT102), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT102), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n717), .A2(new_n726), .A3(new_n927), .A4(new_n672), .ZN(new_n928));
  AND4_X1   g0728(.A1(KEYINPUT103), .A2(new_n926), .A3(new_n728), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT31), .B1(new_n727), .B2(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT103), .B1(new_n930), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n730), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n885), .A2(new_n891), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n914), .A2(new_n852), .A3(new_n916), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT40), .A4(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n932), .A2(new_n934), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n885), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT101), .B1(new_n884), .B2(new_n885), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n932), .ZN(new_n943));
  INV_X1    g0743(.A(new_n442), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n708), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n942), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n863), .B1(new_n925), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n925), .B2(new_n947), .ZN(new_n949));
  INV_X1    g0749(.A(new_n532), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(G116), .A4(new_n215), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n373), .A2(G77), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n240), .B1(new_n211), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n742), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n678), .A2(new_n687), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n636), .A2(new_n562), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n537), .A2(new_n672), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n653), .A2(new_n672), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n959), .A2(KEYINPUT42), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n554), .B1(new_n965), .B2(new_n646), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n673), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT42), .B1(new_n959), .B2(new_n965), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n968), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n469), .A2(new_n672), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n649), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT104), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT104), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n634), .A2(new_n974), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n972), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n970), .A2(new_n971), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n684), .A2(new_n964), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT105), .Z(new_n984));
  INV_X1    g0784(.A(KEYINPUT106), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n981), .A2(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n984), .B(new_n985), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n981), .A2(new_n982), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n691), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT107), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n688), .A2(new_n992), .A3(new_n964), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n992), .B1(new_n688), .B2(new_n964), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n995), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  OR3_X1    g0799(.A1(new_n688), .A2(new_n999), .A3(new_n964), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n688), .B2(new_n964), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n684), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n678), .B(new_n687), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n741), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n996), .A2(new_n998), .A3(new_n685), .A4(new_n1002), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1006), .A3(new_n739), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n990), .B1(new_n1008), .B2(new_n739), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n989), .B1(new_n1009), .B2(new_n745), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n756), .B1(new_n207), .B2(new_n429), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n234), .A2(new_n759), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n746), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT108), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n278), .B1(new_n792), .B2(new_n1015), .C1(new_n420), .C2(new_n795), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n806), .B2(G97), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n784), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n788), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT46), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n788), .B2(new_n579), .ZN(new_n1022));
  INV_X1    g0822(.A(G294), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1020), .B(new_n1022), .C1(new_n1023), .C2(new_n841), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1017), .B1(new_n800), .B2(new_n1018), .C1(KEYINPUT110), .C2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(KEYINPUT110), .B2(new_n1024), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n774), .A2(new_n789), .B1(new_n839), .B2(new_n782), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n806), .A2(G77), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n270), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT111), .Z(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT112), .B(G137), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1019), .A2(G58), .B1(new_n1033), .B2(new_n793), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n202), .B2(new_n795), .C1(new_n375), .C2(new_n841), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n239), .A2(new_n1018), .B1(new_n774), .B2(new_n258), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(G143), .C2(new_n814), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1026), .A2(new_n1028), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT47), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n752), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1038), .A2(KEYINPUT47), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1014), .B1(new_n979), .B2(new_n823), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1010), .A2(new_n1042), .ZN(G387));
  AOI21_X1  g0843(.A(new_n692), .B1(new_n739), .B2(new_n1006), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n739), .B2(new_n1006), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n762), .A2(new_n693), .B1(G107), .B2(new_n207), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n231), .A2(new_n288), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n693), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n256), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n759), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1046), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n746), .B1(new_n1054), .B2(new_n757), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n429), .A2(new_n795), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n270), .B1(new_n792), .B2(new_n258), .C1(new_n788), .C2(new_n326), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n426), .C2(new_n797), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n806), .A2(G97), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n773), .A2(G50), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n814), .A2(G159), .B1(new_n784), .B2(G68), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n788), .A2(new_n1023), .B1(new_n795), .B2(new_n800), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n784), .A2(G303), .B1(G311), .B2(new_n797), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n1015), .B2(new_n774), .C1(new_n775), .C2(new_n782), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT49), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n278), .B1(new_n776), .B2(new_n792), .C1(new_n804), .C2(new_n579), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1062), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1055), .B1(new_n1071), .B2(new_n752), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n678), .B2(new_n823), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT114), .Z(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1006), .B2(new_n745), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1045), .A2(new_n1075), .ZN(G393));
  AND2_X1   g0876(.A1(new_n1008), .A2(new_n691), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n739), .A2(new_n1006), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1004), .A2(new_n745), .A3(new_n1007), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n755), .B(new_n752), .C1(G97), .C2(new_n690), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n238), .A2(new_n759), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n768), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n270), .B1(new_n788), .B2(new_n202), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G143), .B2(new_n793), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n239), .B2(new_n841), .C1(new_n326), .C2(new_n795), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n838), .B(new_n1088), .C1(new_n426), .C2(new_n784), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n774), .A2(new_n375), .B1(new_n258), .B2(new_n782), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n774), .A2(new_n839), .B1(new_n1015), .B2(new_n782), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n278), .B1(new_n788), .B2(new_n800), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G322), .B2(new_n793), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n796), .A2(G116), .B1(G303), .B2(new_n797), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n807), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G294), .B2(new_n784), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1089), .A2(new_n1091), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1085), .B1(new_n820), .B2(new_n1099), .C1(new_n964), .C2(new_n823), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1082), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1081), .A2(new_n1102), .ZN(G390));
  INV_X1    g0903(.A(KEYINPUT115), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n894), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n885), .B2(new_n891), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n701), .A2(new_n700), .B1(new_n637), .B2(new_n704), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n672), .B1(new_n1107), .B2(new_n703), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n918), .B1(new_n1108), .B2(new_n852), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1104), .B(new_n1106), .C1(new_n1109), .C2(new_n917), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n706), .A2(new_n673), .A3(new_n852), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n917), .B1(new_n1111), .B2(new_n919), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n933), .A2(new_n894), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT115), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n893), .B1(new_n920), .B2(new_n1105), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n595), .A2(new_n603), .A3(new_n611), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n666), .A2(new_n675), .A3(new_n477), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1117), .A2(new_n960), .A3(new_n1118), .A4(new_n673), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n727), .A2(new_n728), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n731), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n915), .B1(new_n913), .B2(new_n911), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(G330), .A4(new_n852), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1115), .A2(new_n1116), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n918), .B1(new_n737), .B2(new_n852), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n894), .B1(new_n1125), .B2(new_n917), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n893), .A2(new_n1126), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n932), .A2(G330), .A3(new_n934), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1124), .B(new_n745), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT116), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1124), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n932), .A2(new_n442), .A3(G330), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n626), .B(new_n1133), .C1(new_n922), .C2(new_n944), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1125), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1122), .B1(new_n732), .B2(new_n852), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1123), .A2(new_n919), .A3(new_n1111), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n932), .A2(G330), .A3(new_n852), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n1122), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1134), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1132), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(new_n1124), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n691), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n893), .A2(new_n753), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n746), .B1(new_n828), .B2(new_n426), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n270), .B1(new_n792), .B2(new_n1148), .C1(new_n841), .C2(new_n1032), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G159), .B2(new_n796), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n788), .A2(new_n258), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n239), .C2(new_n804), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G132), .A2(new_n773), .B1(new_n784), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n782), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n270), .B(new_n809), .C1(G294), .C2(new_n793), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n796), .A2(G77), .B1(G107), .B2(new_n797), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n834), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G97), .A2(new_n784), .B1(new_n773), .B2(G116), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n800), .B2(new_n782), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1153), .A2(new_n1158), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1147), .B1(new_n1164), .B2(new_n752), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1146), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1131), .A2(new_n1145), .A3(new_n1166), .ZN(G378));
  NAND2_X1  g0967(.A1(new_n940), .A2(new_n941), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n267), .A2(new_n670), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n316), .B(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1168), .A2(new_n1173), .A3(G330), .A4(new_n935), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n932), .A2(new_n934), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n904), .B2(new_n905), .ZN(new_n1176));
  OAI211_X1 g0976(.A(G330), .B(new_n935), .C1(new_n1176), .C2(KEYINPUT40), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1172), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1174), .A2(new_n1178), .A3(new_n921), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n921), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n745), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1172), .A2(new_n753), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n746), .B1(new_n828), .B2(G50), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n239), .B1(G33), .B2(G41), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n278), .B2(new_n287), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n420), .A2(new_n774), .B1(new_n1018), .B2(new_n429), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G116), .B2(new_n814), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n806), .A2(G58), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n841), .A2(new_n460), .B1(new_n795), .B2(new_n202), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n788), .A2(new_n326), .B1(new_n800), .B2(new_n792), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1189), .A2(new_n1190), .A3(G41), .A4(new_n270), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1019), .A2(new_n1155), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n796), .A2(G150), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n797), .A2(G132), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n774), .A2(new_n1157), .B1(new_n1148), .B2(new_n782), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G137), .C2(new_n784), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT59), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1195), .B1(new_n375), .B2(new_n804), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1201), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1194), .B1(new_n1193), .B2(new_n1192), .C1(new_n1203), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1183), .B1(new_n1206), .B2(new_n752), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1182), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1181), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n921), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1173), .B1(new_n942), .B2(G330), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1177), .A2(new_n1172), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1174), .A2(new_n1178), .A3(new_n921), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1210), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1134), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1144), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n692), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1218), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1210), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1209), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G375));
  NOR2_X1   g1023(.A1(new_n1141), .A2(new_n990), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1137), .A2(new_n1140), .A3(new_n1134), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n745), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n768), .B1(new_n827), .B2(new_n202), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1056), .B1(new_n773), .B2(G283), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT117), .Z(new_n1231));
  OAI221_X1 g1031(.A(new_n278), .B1(new_n792), .B2(new_n789), .C1(new_n788), .C2(new_n460), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G116), .B2(new_n797), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n814), .A2(G294), .B1(new_n784), .B2(G107), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1231), .A2(new_n1029), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n814), .A2(G132), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT118), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n270), .B1(new_n788), .B2(new_n375), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n841), .A2(new_n1154), .B1(new_n239), .B2(new_n795), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G128), .C2(new_n793), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G150), .A2(new_n784), .B1(new_n773), .B2(new_n1033), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1237), .A2(new_n1188), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT119), .B1(new_n1235), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1235), .A2(KEYINPUT119), .A3(new_n1242), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n752), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1229), .B1(new_n1243), .B2(new_n1245), .C1(new_n1122), .C2(new_n754), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1228), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1226), .A2(new_n1248), .ZN(G381));
  NOR2_X1   g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1226), .A2(new_n1248), .A3(new_n861), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(G387), .A2(G390), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT120), .Z(new_n1254));
  INV_X1    g1054(.A(G378), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1222), .A2(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1254), .A2(new_n1256), .ZN(G407));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1247), .B1(new_n861), .B2(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1225), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT60), .B1(new_n1225), .B2(KEYINPUT123), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n691), .B(new_n1142), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n861), .A2(new_n1260), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1267), .A2(new_n1268), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1275), .A2(new_n745), .B1(new_n1182), .B2(new_n1207), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT122), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT122), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1209), .A2(new_n1278), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1220), .A2(new_n990), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1255), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT121), .B1(new_n1222), .B2(G378), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1218), .B(KEYINPUT57), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1214), .A2(new_n1215), .B1(new_n1217), .B2(new_n1144), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1284), .B(new_n691), .C1(new_n1285), .C2(KEYINPUT57), .ZN(new_n1286));
  AND4_X1   g1086(.A1(KEYINPUT121), .A2(new_n1286), .A3(G378), .A4(new_n1276), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1282), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n671), .A2(G213), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1274), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1259), .B1(new_n1290), .B2(KEYINPUT61), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1286), .A2(G378), .A3(new_n1276), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT121), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1222), .A2(KEYINPUT121), .A3(G378), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1297), .A2(new_n1282), .B1(G213), .B2(new_n671), .ZN(new_n1298));
  OAI211_X1 g1098(.A(KEYINPUT127), .B(new_n1292), .C1(new_n1298), .C2(new_n1274), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1288), .A2(new_n1289), .A3(new_n1269), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1298), .A2(new_n1302), .A3(new_n1269), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1291), .A2(new_n1299), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1101), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G387), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G390), .A2(new_n1010), .A3(new_n1042), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT126), .B1(G387), .B2(new_n1305), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n825), .B1(new_n1045), .B2(new_n1075), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1250), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1308), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1306), .A2(new_n1307), .A3(KEYINPUT126), .A4(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1304), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1274), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1318), .B2(new_n1317), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1269), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1300), .A2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1315), .A2(KEYINPUT61), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(new_n1321), .A3(new_n1323), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(G405));
  AOI22_X1  g1126(.A1(new_n1295), .A2(new_n1296), .B1(new_n1255), .B2(G375), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1315), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1315), .A2(new_n1327), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1328), .A2(new_n1329), .B1(new_n1268), .B2(new_n1267), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1315), .A2(new_n1327), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1315), .A2(new_n1327), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1269), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1330), .A2(new_n1333), .ZN(G402));
endmodule


