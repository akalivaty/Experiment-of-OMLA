//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368, new_n1369, new_n1370;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT66), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n207), .B2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G13), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n221), .A2(KEYINPUT66), .A3(G1), .A4(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(new_n209), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n218), .A2(new_n225), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G232), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G107), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n260), .A2(new_n210), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n248), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n268), .A3(G274), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n265), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(KEYINPUT67), .A3(new_n265), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G244), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n263), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n230), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n229), .A2(new_n256), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n281), .A2(new_n282), .B1(new_n229), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT15), .B(G87), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n229), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n280), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n280), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(G77), .B1(new_n229), .B2(G1), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n288), .B1(G77), .B2(new_n289), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n278), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n276), .A2(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(new_n276), .B2(G200), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n263), .A2(G190), .A3(new_n269), .A4(new_n275), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT69), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n274), .A2(G226), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n269), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n252), .A2(G222), .B1(G77), .B2(new_n251), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT68), .B(G223), .Z(new_n308));
  OR2_X1    g0108(.A1(new_n260), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n268), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n306), .A2(new_n310), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G190), .ZN(new_n314));
  INV_X1    g0114(.A(new_n280), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT8), .B(G58), .Z(new_n316));
  INV_X1    g0116(.A(new_n286), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G20), .A2(G33), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n316), .A2(new_n317), .B1(G150), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n203), .A2(G20), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G50), .B1(new_n229), .B2(G1), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n292), .A2(new_n322), .B1(G50), .B2(new_n289), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n324), .A2(KEYINPUT9), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(KEYINPUT9), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n312), .A2(new_n314), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT10), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(new_n314), .A4(new_n312), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n311), .A2(new_n277), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n313), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n324), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n304), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n281), .B1(new_n264), .B2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n291), .B1(new_n290), .B2(new_n281), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n251), .B2(new_n229), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n258), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G58), .A2(G68), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n346), .B2(new_n202), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT75), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n318), .A2(G159), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n229), .B1(new_n227), .B2(new_n345), .ZN(new_n351));
  INV_X1    g0151(.A(G159), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n282), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT75), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n344), .A2(KEYINPUT16), .A3(new_n350), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n280), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n257), .A2(new_n229), .A3(new_n258), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n342), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n343), .A2(KEYINPUT76), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(G68), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n354), .A2(new_n350), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT16), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n340), .B1(new_n356), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G226), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G1698), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n368), .B1(G223), .B2(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n248), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n268), .A2(G232), .A3(new_n265), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n269), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n277), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n268), .B1(new_n369), .B2(new_n370), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n377), .A2(new_n374), .A3(new_n334), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n366), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n366), .A2(new_n383), .A3(new_n380), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n372), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G200), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n377), .B2(new_n374), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n340), .B(new_n389), .C1(new_n356), .C2(new_n365), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n363), .A2(new_n364), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n354), .A2(new_n350), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n209), .B1(new_n359), .B2(new_n342), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n315), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n340), .A4(new_n389), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n382), .A2(new_n384), .A3(new_n392), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT11), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n209), .A2(G20), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n286), .B2(new_n283), .ZN(new_n405));
  INV_X1    g0205(.A(G50), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT71), .B1(new_n282), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n318), .A2(new_n408), .A3(G50), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n403), .B1(new_n410), .B2(new_n315), .ZN(new_n411));
  INV_X1    g0211(.A(new_n409), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n408), .B1(new_n318), .B2(G50), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT11), .B(new_n280), .C1(new_n414), .C2(new_n405), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT12), .B1(new_n289), .B2(G68), .ZN(new_n416));
  OR3_X1    g0216(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n209), .B1(new_n264), .B2(G20), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n416), .A2(new_n417), .B1(new_n291), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n411), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT72), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT72), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n411), .A2(new_n415), .A3(new_n422), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(G226), .A2(G1698), .ZN(new_n425));
  INV_X1    g0225(.A(G232), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G1698), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n259), .B1(G33), .B2(G97), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n269), .B1(new_n428), .B2(new_n268), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n210), .B1(new_n272), .B2(new_n273), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT13), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G226), .B2(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G97), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n433), .A2(new_n251), .B1(new_n256), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G274), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n248), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n435), .A2(new_n248), .B1(new_n437), .B2(new_n266), .ZN(new_n438));
  INV_X1    g0238(.A(new_n273), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT67), .B1(new_n268), .B2(new_n265), .ZN(new_n440));
  OAI21_X1  g0240(.A(G238), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n277), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT70), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n442), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n429), .B2(new_n430), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n438), .A2(new_n448), .A3(new_n441), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n444), .A2(new_n445), .B1(new_n452), .B2(G179), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n424), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n429), .A2(new_n430), .A3(new_n449), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n448), .B1(new_n438), .B2(new_n441), .ZN(new_n457));
  OAI21_X1  g0257(.A(G190), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT13), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n442), .B1(new_n438), .B2(new_n441), .ZN(new_n460));
  OAI21_X1  g0260(.A(G200), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n424), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT73), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n424), .A2(new_n458), .A3(new_n461), .A4(KEYINPUT73), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n455), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n338), .A2(new_n402), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT5), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n264), .B(G45), .C1(new_n470), .C2(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(KEYINPUT79), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G257), .B(new_n268), .C1(new_n473), .C2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n474), .A3(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(KEYINPUT79), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n437), .A2(new_n481), .A3(new_n482), .A4(new_n471), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G1698), .ZN(new_n485));
  OAI211_X1 g0285(.A(G244), .B(new_n485), .C1(new_n249), .C2(new_n250), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n248), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n484), .A2(new_n334), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n480), .A2(new_n483), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n248), .B2(new_n492), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(G169), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n361), .A2(G107), .A3(new_n362), .ZN(new_n498));
  XOR2_X1   g0298(.A(G97), .B(G107), .Z(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT77), .B(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n261), .A2(KEYINPUT6), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n499), .A2(KEYINPUT6), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G20), .B1(G77), .B2(new_n318), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n315), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n289), .A2(G97), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT78), .B1(new_n256), .B2(G1), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n264), .A3(G33), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n291), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n506), .B1(new_n511), .B2(new_n434), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n469), .B1(new_n497), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n504), .A2(new_n512), .ZN(new_n515));
  AOI21_X1  g0315(.A(G169), .B1(new_n484), .B2(new_n493), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n515), .A2(KEYINPUT80), .A3(new_n494), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n484), .A2(new_n493), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G200), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n513), .B(new_n520), .C1(new_n385), .C2(new_n519), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n514), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n523));
  OAI211_X1 g0323(.A(G250), .B(new_n485), .C1(new_n249), .C2(new_n250), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n256), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n248), .ZN(new_n527));
  OAI211_X1 g0327(.A(G264), .B(new_n268), .C1(new_n473), .C2(new_n479), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n483), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n387), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n527), .A2(new_n385), .A3(new_n483), .A4(new_n528), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n229), .B1(new_n249), .B2(new_n250), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G87), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n536), .ZN(new_n538));
  INV_X1    g0338(.A(new_n533), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n259), .A2(new_n538), .A3(new_n229), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n229), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n261), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT81), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n229), .A3(G33), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n537), .A2(new_n540), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT24), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n256), .B1(new_n546), .B2(new_n548), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n229), .B1(new_n542), .B2(new_n543), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n540), .A4(new_n537), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n280), .ZN(new_n558));
  INV_X1    g0358(.A(new_n511), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n289), .A2(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT25), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n532), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n527), .A2(new_n334), .A3(new_n483), .A4(new_n528), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n529), .A2(new_n277), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n315), .B1(new_n552), .B2(new_n556), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n563), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n212), .B1(new_n475), .B2(G1), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n264), .A2(new_n436), .A3(G45), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n268), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n547), .A2(G116), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n545), .A2(KEYINPUT81), .ZN(new_n574));
  OAI21_X1  g0374(.A(G33), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n576));
  OAI211_X1 g0376(.A(G238), .B(new_n485), .C1(new_n249), .C2(new_n250), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n578), .B2(new_n248), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n277), .ZN(new_n580));
  AOI211_X1 g0380(.A(new_n334), .B(new_n572), .C1(new_n578), .C2(new_n248), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT82), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n248), .ZN(new_n583));
  INV_X1    g0383(.A(new_n572), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(G179), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n277), .C2(new_n579), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n500), .B2(new_n286), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n259), .A2(new_n229), .A3(G68), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G87), .A2(G107), .ZN(new_n592));
  NAND3_X1  g0392(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n500), .A2(new_n592), .B1(new_n229), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n280), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n285), .A2(new_n290), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n511), .C2(new_n285), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n582), .A2(new_n587), .A3(new_n597), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n385), .B(new_n572), .C1(new_n578), .C2(new_n248), .ZN(new_n599));
  INV_X1    g0399(.A(new_n579), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(G200), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n559), .A2(G87), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(new_n602), .A3(new_n596), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n565), .A2(new_n569), .A3(new_n598), .A4(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n510), .A2(new_n315), .A3(G116), .A4(new_n289), .ZN(new_n607));
  XNOR2_X1  g0407(.A(KEYINPUT81), .B(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n290), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT20), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n280), .B1(new_n549), .B2(new_n229), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n490), .A2(new_n229), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n434), .A2(KEYINPUT77), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT77), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G97), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n617), .B2(new_n256), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n611), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n229), .B(new_n490), .C1(new_n500), .C2(G33), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n608), .A2(G20), .B1(new_n230), .B2(new_n279), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT20), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n610), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n624));
  OAI211_X1 g0424(.A(G257), .B(new_n485), .C1(new_n249), .C2(new_n250), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n257), .A2(G303), .A3(new_n258), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n248), .ZN(new_n628));
  OAI211_X1 g0428(.A(G270), .B(new_n268), .C1(new_n473), .C2(new_n479), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n483), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n623), .A2(new_n630), .A3(new_n334), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(G200), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n633), .B(new_n623), .C1(new_n385), .C2(new_n630), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n607), .A2(new_n609), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n612), .A2(new_n618), .A3(new_n611), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT20), .B1(new_n620), .B2(new_n621), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n639));
  AND4_X1   g0439(.A1(G169), .A2(new_n638), .A3(new_n630), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n619), .A2(new_n622), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n277), .B1(new_n641), .B2(new_n635), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n630), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n632), .B(new_n634), .C1(new_n640), .C2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n606), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n468), .A2(new_n522), .A3(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n337), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n366), .A2(new_n383), .A3(new_n380), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n383), .B1(new_n366), .B2(new_n380), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n295), .A2(new_n296), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n454), .B1(new_n651), .B2(new_n462), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n390), .B(KEYINPUT17), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n647), .B1(new_n655), .B2(new_n332), .ZN(new_n656));
  INV_X1    g0456(.A(new_n468), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n585), .B1(new_n277), .B2(new_n579), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n597), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n601), .A2(new_n604), .B1(new_n658), .B2(new_n597), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n565), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n638), .A2(G169), .A3(new_n630), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(KEYINPUT83), .B2(KEYINPUT21), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n642), .A2(new_n630), .A3(new_n639), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n631), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n662), .B1(new_n666), .B2(new_n569), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n660), .B1(new_n667), .B2(new_n522), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n484), .A2(new_n334), .A3(new_n493), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n516), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n661), .A2(new_n669), .A3(new_n671), .A4(new_n515), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n598), .A2(new_n605), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT80), .B1(new_n671), .B2(new_n515), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n497), .A2(new_n469), .A3(new_n513), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n673), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n668), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n656), .B1(new_n657), .B2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n264), .A2(new_n229), .A3(G13), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n682), .A2(KEYINPUT85), .A3(KEYINPUT27), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT85), .B1(new_n682), .B2(KEYINPUT27), .ZN(new_n684));
  OAI221_X1 g0484(.A(G213), .B1(KEYINPUT27), .B2(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n666), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n565), .A2(new_n569), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n569), .B2(new_n687), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT86), .Z(new_n692));
  INV_X1    g0492(.A(new_n666), .ZN(new_n693));
  INV_X1    g0493(.A(new_n687), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n623), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n644), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n687), .B1(new_n568), .B2(new_n563), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n689), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n569), .B2(new_n694), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n692), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT87), .Z(G399));
  INV_X1    g0505(.A(new_n223), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n706), .A2(KEYINPUT88), .A3(G41), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT88), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n223), .B2(new_n470), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n500), .A2(new_n545), .A3(new_n592), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n264), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n228), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n710), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  NAND2_X1  g0515(.A1(new_n671), .A2(new_n515), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n605), .A2(new_n659), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n716), .A2(new_n717), .A3(new_n669), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n677), .B2(new_n669), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n661), .A2(new_n565), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n569), .B(new_n632), .C1(new_n643), .C2(new_n640), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n514), .A2(new_n518), .A3(new_n521), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n659), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n694), .C1(new_n719), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n687), .B1(new_n668), .B2(new_n678), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(KEYINPUT29), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n723), .A2(new_n606), .A3(new_n644), .A4(new_n687), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n628), .A2(new_n629), .A3(new_n483), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n493), .A3(new_n484), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n581), .A2(new_n528), .A3(new_n527), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n527), .A2(new_n528), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n585), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n496), .A3(KEYINPUT30), .A4(new_n730), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n579), .A2(G179), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n519), .A2(new_n630), .A3(new_n529), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n687), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(G330), .B1(new_n728), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n727), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n715), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n710), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n221), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n264), .B1(new_n749), .B2(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OR3_X1    g0551(.A1(KEYINPUT91), .A2(G13), .A3(G33), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT91), .B1(G13), .B2(G33), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n230), .B1(G20), .B2(new_n277), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n243), .A2(new_n475), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n223), .A2(new_n251), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT89), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n475), .B2(new_n713), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT90), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n706), .A2(new_n251), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n768), .A2(G355), .B1(new_n545), .B2(new_n706), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n759), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n229), .A2(new_n334), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n385), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G326), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n772), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(KEYINPUT33), .A2(G317), .ZN(new_n779));
  NAND2_X1  g0579(.A1(KEYINPUT33), .A2(G317), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n385), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n229), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n776), .B(new_n781), .C1(G294), .C2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n771), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n385), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n229), .A2(G190), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(new_n334), .A3(new_n387), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n787), .A2(G322), .B1(G329), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n791), .B(new_n251), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n334), .A2(G200), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT92), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n797), .A2(new_n229), .A3(G190), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(G283), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n797), .A2(new_n229), .A3(new_n385), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n785), .B(new_n799), .C1(new_n800), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n783), .A2(new_n434), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n790), .A2(G159), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n809), .B2(KEYINPUT32), .C1(new_n209), .C2(new_n778), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n798), .A2(G107), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n802), .B2(new_n211), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n809), .A2(KEYINPUT32), .B1(G50), .B2(new_n773), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n251), .B1(new_n793), .B2(G77), .ZN(new_n814));
  INV_X1    g0614(.A(new_n787), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n814), .C1(new_n226), .C2(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n806), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n751), .B(new_n770), .C1(new_n757), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n756), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n697), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n697), .A2(G330), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n698), .A2(new_n751), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(G396));
  INV_X1    g0624(.A(new_n751), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n297), .A2(new_n303), .A3(new_n694), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n598), .A2(new_n605), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n514), .B2(new_n518), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n672), .B1(new_n828), .B2(new_n669), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n724), .B2(new_n829), .ZN(new_n830));
  AND4_X1   g0630(.A1(new_n294), .A2(new_n296), .A3(new_n278), .A4(new_n694), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n294), .A2(new_n687), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n303), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n297), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n726), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n825), .B1(new_n835), .B2(new_n745), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n745), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n757), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n755), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n825), .B1(G77), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n805), .A2(new_n261), .ZN(new_n842));
  INV_X1    g0642(.A(new_n798), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n211), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n251), .B1(new_n789), .B2(new_n792), .C1(new_n815), .C2(new_n525), .ZN(new_n845));
  NOR4_X1   g0645(.A1(new_n842), .A2(new_n807), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n549), .A2(new_n793), .B1(new_n773), .B2(G303), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n778), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT94), .Z(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n787), .B1(new_n793), .B2(G159), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n777), .A2(G150), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n774), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n855));
  XNOR2_X1  g0655(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n798), .A2(G68), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n251), .B1(new_n790), .B2(G132), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n226), .C2(new_n783), .ZN(new_n859));
  INV_X1    g0659(.A(new_n805), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(G50), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n846), .A2(new_n850), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n841), .B1(new_n834), .B2(new_n755), .C1(new_n838), .C2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n837), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n749), .A2(new_n264), .ZN(new_n866));
  INV_X1    g0666(.A(G330), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n728), .A2(new_n744), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n424), .A2(new_n694), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n444), .A2(new_n445), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n452), .A2(G179), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n444), .A2(new_n445), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n870), .B1(new_n466), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n462), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n454), .A2(new_n877), .A3(new_n869), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n834), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n868), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n340), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n395), .B2(new_n399), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n390), .B1(new_n883), .B2(new_n379), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n685), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT99), .ZN(new_n887));
  INV_X1    g0687(.A(new_n685), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n366), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n381), .A2(new_n889), .A3(new_n890), .A4(new_n390), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n887), .B1(new_n886), .B2(new_n891), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n401), .A2(new_n392), .A3(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n382), .A3(new_n384), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT100), .B1(new_n401), .B2(new_n392), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n885), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n355), .A3(new_n280), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n685), .B1(new_n902), .B2(new_n340), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n650), .B2(new_n653), .ZN(new_n905));
  INV_X1    g0705(.A(new_n390), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n340), .A2(new_n902), .B1(new_n379), .B2(new_n685), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n891), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n881), .B(KEYINPUT101), .C1(new_n900), .C2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n886), .A2(new_n891), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT99), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n899), .A2(new_n915), .A3(new_n892), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n911), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n295), .A2(new_n296), .A3(new_n694), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n299), .B(new_n300), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n298), .B1(new_n294), .B2(new_n687), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n920), .B2(new_n651), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n431), .A2(new_n443), .ZN(new_n922));
  AOI22_X1  g0722(.A1(G190), .A2(new_n452), .B1(new_n922), .B2(G200), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT73), .B1(new_n923), .B2(new_n424), .ZN(new_n924));
  INV_X1    g0724(.A(new_n465), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n875), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n869), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n455), .A2(new_n462), .A3(new_n870), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n921), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n645), .A2(new_n522), .A3(new_n694), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT31), .B1(new_n739), .B2(new_n687), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(KEYINPUT40), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n913), .B1(new_n917), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n910), .B1(new_n905), .B2(new_n909), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n402), .A2(new_n903), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n891), .A2(new_n908), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(KEYINPUT38), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n934), .A3(new_n929), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n912), .A2(new_n936), .B1(new_n880), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n657), .A2(new_n868), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n867), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT102), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n830), .A2(new_n918), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n876), .A2(new_n878), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n685), .B1(new_n648), .B2(new_n649), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT98), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(KEYINPUT98), .A3(new_n953), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n937), .B2(new_n940), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n916), .A2(new_n910), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n940), .A2(new_n957), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n454), .A2(new_n694), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n955), .A2(new_n956), .A3(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n468), .B(new_n725), .C1(new_n726), .C2(KEYINPUT29), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n656), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n866), .B1(new_n948), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n948), .B2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n713), .A2(G77), .A3(new_n345), .ZN(new_n973));
  INV_X1    g0773(.A(new_n201), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n209), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(G1), .A3(new_n221), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n230), .A2(new_n229), .A3(new_n545), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT96), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n972), .A2(new_n976), .A3(new_n984), .ZN(G367));
  INV_X1    g0785(.A(new_n703), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n522), .B1(new_n513), .B2(new_n694), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n716), .B2(new_n694), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT104), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n603), .A2(new_n687), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT103), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n659), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n661), .B2(new_n992), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n990), .B(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n994), .A2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n690), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n988), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT42), .Z(new_n1001));
  INV_X1    g0801(.A(new_n569), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n988), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n514), .A2(new_n518), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n694), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n998), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n997), .B(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n710), .B(KEYINPUT41), .Z(new_n1008));
  OR2_X1    g0808(.A1(new_n692), .A2(new_n988), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n692), .A2(new_n988), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT105), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT105), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n692), .A2(new_n1014), .A3(new_n988), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1011), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n986), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n702), .A2(new_n688), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n999), .B1(new_n1022), .B2(KEYINPUT106), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(KEYINPUT106), .B2(new_n1022), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(new_n699), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1011), .A2(new_n1019), .A3(new_n703), .A4(new_n1016), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1021), .A2(new_n746), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1008), .B1(new_n1027), .B2(new_n746), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n750), .B(KEYINPUT107), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n1007), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n763), .A2(new_n239), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n758), .B1(new_n223), .B2(new_n285), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n825), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n805), .A2(new_n1034), .A3(new_n545), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n787), .A2(G303), .B1(G317), .B2(new_n790), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n251), .C1(new_n848), .C2(new_n794), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n617), .B2(new_n798), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1034), .B1(new_n802), .B2(new_n608), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n774), .A2(new_n792), .B1(new_n261), .B2(new_n783), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G294), .B2(new_n777), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n974), .A2(new_n793), .B1(new_n787), .B2(G150), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n853), .B2(new_n789), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G58), .B2(new_n801), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n259), .B1(new_n843), .B2(new_n283), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT108), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n783), .A2(new_n209), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n352), .B2(new_n778), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G143), .B2(new_n773), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1045), .A2(new_n1048), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1035), .A2(new_n1042), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT47), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1033), .B1(new_n1056), .B2(new_n757), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n994), .A2(new_n756), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1030), .A2(new_n1059), .ZN(G387));
  OR2_X1    g0860(.A1(new_n702), .A2(new_n820), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n762), .B1(new_n236), .B2(new_n475), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n711), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n768), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n281), .A2(G50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g0867(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1065), .A2(new_n1069), .B1(new_n261), .B2(new_n706), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n825), .B1(new_n1070), .B2(new_n759), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G303), .A2(new_n793), .B1(new_n787), .B2(G317), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n773), .A2(G322), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n792), .C2(new_n778), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT48), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n801), .A2(G294), .B1(G283), .B2(new_n784), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT109), .Z(new_n1077));
  NOR2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(KEYINPUT49), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n251), .B1(new_n789), .B2(new_n775), .C1(new_n843), .C2(new_n608), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(KEYINPUT49), .B2(new_n1078), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n783), .A2(new_n285), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G159), .B2(new_n773), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n281), .B2(new_n778), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n801), .A2(G77), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n251), .B1(new_n793), .B2(G68), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n787), .A2(G50), .B1(G150), .B2(new_n790), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n434), .B2(new_n843), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1082), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1071), .B1(new_n1091), .B2(new_n757), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1025), .A2(new_n1029), .B1(new_n1061), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1025), .A2(new_n746), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n710), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1025), .A2(new_n746), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(new_n1021), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1026), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n710), .A3(new_n1027), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT110), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT110), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1021), .A2(new_n1103), .A3(new_n1026), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1029), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n763), .A2(new_n246), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n758), .B1(new_n223), .B2(new_n500), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n825), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n783), .A2(new_n283), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n790), .A2(G143), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n259), .B(new_n1110), .C1(new_n794), .C2(new_n281), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n974), .C2(new_n777), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n209), .B2(new_n802), .C1(new_n211), .C2(new_n843), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n787), .A2(G159), .B1(new_n773), .B2(G150), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT51), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n778), .A2(new_n800), .B1(new_n608), .B2(new_n783), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n251), .B1(new_n794), .B2(new_n525), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G322), .C2(new_n790), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n811), .C1(new_n848), .C2(new_n802), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n787), .A2(G311), .B1(new_n773), .B2(G317), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1113), .A2(new_n1115), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT112), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n838), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1108), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n988), .B2(new_n820), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1101), .A2(new_n1105), .A3(new_n1128), .ZN(G390));
  AOI21_X1  g0929(.A(new_n831), .B1(new_n679), .B2(new_n826), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n964), .B1(new_n1130), .B2(new_n950), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n962), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n833), .A2(new_n297), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n694), .B(new_n1133), .C1(new_n719), .C2(new_n724), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n918), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n951), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n959), .A2(new_n940), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n964), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n867), .B1(new_n930), .B2(new_n933), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n929), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1132), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT113), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1139), .A2(new_n929), .A3(KEYINPUT113), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1029), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n825), .B1(new_n316), .B2(new_n839), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n787), .A2(G132), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n259), .B1(new_n794), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(G125), .C2(new_n790), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n778), .A2(new_n853), .B1(new_n352), .B2(new_n783), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G128), .B2(new_n773), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(new_n201), .C2(new_n843), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n801), .A2(G150), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT53), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n805), .A2(new_n211), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n774), .A2(new_n848), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1109), .B(new_n1160), .C1(G107), .C2(new_n777), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n259), .B1(new_n790), .B2(G294), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n617), .A2(new_n793), .B1(new_n787), .B2(G116), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1161), .A2(new_n857), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1156), .A2(new_n1158), .B1(new_n1159), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1149), .B1(new_n1165), .B2(new_n757), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n963), .B2(new_n755), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n968), .B(new_n656), .C1(new_n657), .C2(new_n745), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n950), .B1(new_n745), .B2(new_n921), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n745), .A2(new_n879), .A3(new_n1142), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT113), .B1(new_n1139), .B2(new_n929), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n949), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT114), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n834), .B1(new_n745), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1139), .A2(KEYINPUT114), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n950), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1140), .A2(new_n918), .A3(new_n1134), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1168), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT116), .B1(new_n1147), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1132), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n917), .A2(new_n965), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1136), .A2(new_n1183), .B1(new_n962), .B2(new_n1131), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1184), .B2(new_n1145), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT116), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1168), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1130), .B1(new_n1145), .B2(new_n1169), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1140), .A2(new_n918), .A3(new_n1134), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n921), .B1(new_n1139), .B2(KEYINPUT114), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(KEYINPUT114), .B2(new_n1139), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n1191), .B2(new_n950), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1187), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1185), .A2(new_n1186), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n748), .B1(new_n1181), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT117), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT115), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1145), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n965), .B1(new_n949), .B2(new_n951), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n960), .B1(new_n910), .B2(new_n916), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1199), .A2(new_n958), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n950), .B1(new_n1134), .B2(new_n918), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1202), .A2(new_n917), .A3(new_n965), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1198), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT115), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1180), .A2(new_n1204), .A3(new_n1205), .A4(new_n1182), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1197), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1195), .A2(new_n1196), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1196), .B1(new_n1195), .B2(new_n1207), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1148), .B(new_n1167), .C1(new_n1208), .C2(new_n1209), .ZN(G378));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n1147), .B2(new_n1180), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1205), .A2(new_n1180), .A3(new_n1204), .A4(new_n1182), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1187), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n912), .A2(new_n936), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n867), .B1(new_n942), .B2(new_n880), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT120), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(KEYINPUT120), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n332), .A2(new_n337), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n336), .A2(new_n888), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT55), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1220), .B(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1224));
  XOR2_X1   g1024(.A(new_n1223), .B(new_n1224), .Z(new_n1225));
  NAND3_X1  g1025(.A1(new_n1218), .A2(new_n1219), .A3(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n955), .A2(new_n956), .A3(new_n966), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1225), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1228), .A2(KEYINPUT120), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1214), .A2(new_n1215), .A3(KEYINPUT120), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT120), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1228), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1229), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n967), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1230), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT121), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1230), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1168), .B1(new_n1197), .B2(new_n1206), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1226), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1227), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT121), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1238), .B1(new_n1207), .B2(new_n1187), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1237), .A2(new_n710), .A3(new_n1241), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1228), .A2(new_n754), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n825), .B1(new_n974), .B2(new_n839), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1050), .B1(new_n545), .B2(new_n774), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n798), .A2(G58), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n251), .A2(new_n470), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n285), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n793), .B2(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n787), .A2(G107), .B1(G283), .B2(new_n790), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1086), .A2(new_n1252), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1251), .B(new_n1257), .C1(G97), .C2(new_n777), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT58), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1253), .B(new_n406), .C1(G33), .C2(G41), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT118), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n787), .A2(G128), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n794), .B2(new_n853), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G132), .B2(new_n777), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G150), .A2(new_n784), .B1(new_n773), .B2(G125), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n802), .C2(new_n1151), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(KEYINPUT59), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(KEYINPUT59), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n798), .A2(G159), .ZN(new_n1270));
  AOI211_X1 g1070(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1262), .B1(KEYINPUT58), .B2(new_n1258), .C1(new_n1268), .C2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1250), .B1(new_n1273), .B2(new_n757), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1244), .A2(new_n1029), .B1(new_n1249), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1248), .A2(new_n1275), .ZN(G375));
  OAI21_X1  g1076(.A(new_n1029), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT122), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n825), .B1(G68), .B2(new_n839), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n778), .A2(new_n1151), .B1(new_n406), .B2(new_n783), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G132), .B2(new_n773), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n251), .B1(new_n790), .B2(G128), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G137), .A2(new_n787), .B1(new_n793), .B2(G150), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1252), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1281), .B(new_n1284), .C1(new_n805), .C2(new_n352), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n251), .B1(new_n789), .B2(new_n800), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n525), .A2(new_n774), .B1(new_n778), .B2(new_n608), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1286), .B(new_n1287), .C1(G107), .C2(new_n793), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1083), .B1(G283), .B2(new_n787), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(KEYINPUT123), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1288), .B(new_n1290), .C1(new_n283), .C2(new_n843), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n805), .A2(new_n434), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1279), .B1(new_n1293), .B2(new_n757), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n951), .B2(new_n755), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(KEYINPUT122), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1278), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1180), .A2(new_n1008), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1168), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1298), .A2(new_n1302), .ZN(G381));
  INV_X1    g1103(.A(G390), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1298), .A3(new_n1302), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1148), .A2(new_n1167), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1195), .B2(new_n1207), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  OR4_X1    g1109(.A1(G387), .A2(new_n1306), .A3(G375), .A4(new_n1309), .ZN(G407));
  NAND2_X1  g1110(.A1(new_n686), .A2(G213), .ZN(new_n1311));
  OR3_X1    g1111(.A1(G375), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G407), .A2(G213), .A3(new_n1312), .ZN(G409));
  NAND3_X1  g1113(.A1(new_n1248), .A2(G378), .A3(new_n1275), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1275), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1239), .A2(new_n1008), .A3(new_n1240), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1308), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1311), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1300), .A2(KEYINPUT60), .A3(new_n1168), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n710), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1193), .A2(KEYINPUT60), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1301), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n864), .B1(new_n1323), .B2(new_n1297), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1323), .A2(new_n864), .A3(new_n1297), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n686), .A2(G213), .A3(G2897), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1327), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT125), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1326), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(new_n1328), .A3(new_n1324), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1334), .A2(G213), .A3(new_n686), .A4(G2897), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1330), .B1(new_n1332), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1336), .ZN(new_n1337));
  OR2_X1    g1137(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1318), .A2(new_n1311), .A3(new_n1327), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  AOI22_X1  g1141(.A1(new_n1314), .A2(new_n1317), .B1(G213), .B2(new_n686), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1338), .B1(new_n1342), .B2(new_n1327), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1337), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT127), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G390), .B1(new_n1030), .B2(new_n1059), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  XOR2_X1   g1147(.A(G393), .B(G396), .Z(new_n1348));
  NAND3_X1  g1148(.A1(G390), .A2(new_n1030), .A3(new_n1059), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1347), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1348), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1349), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1351), .B1(new_n1352), .B2(new_n1346), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1350), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT127), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1355), .B(new_n1337), .C1(new_n1341), .C2(new_n1343), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1345), .A2(new_n1354), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1342), .A2(new_n1327), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1354), .B1(KEYINPUT63), .B2(new_n1359), .ZN(new_n1360));
  NOR3_X1   g1160(.A1(new_n1359), .A2(KEYINPUT124), .A3(KEYINPUT63), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT124), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1362), .B1(new_n1358), .B2(new_n1363), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1360), .B(new_n1337), .C1(new_n1361), .C2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1357), .A2(new_n1365), .ZN(G405));
  INV_X1    g1166(.A(new_n1314), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1309), .B1(new_n1248), .B2(new_n1275), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  XNOR2_X1  g1169(.A(new_n1369), .B(new_n1331), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1370), .B(new_n1354), .ZN(G402));
endmodule


