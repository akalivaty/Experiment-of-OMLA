

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n712), .A2(n711), .ZN(n761) );
  AND2_X1 U556 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U557 ( .A1(n677), .A2(n676), .ZN(n678) );
  BUF_X1 U558 ( .A(n715), .Z(n716) );
  INV_X1 U559 ( .A(G2105), .ZN(n524) );
  NOR2_X2 U560 ( .A1(n534), .A2(n533), .ZN(G160) );
  OR2_X1 U561 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U562 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U563 ( .A(KEYINPUT98), .B(KEYINPUT32), .ZN(n682) );
  XOR2_X1 U564 ( .A(KEYINPUT27), .B(n605), .Z(n523) );
  INV_X1 U565 ( .A(n666), .ZN(n646) );
  INV_X1 U566 ( .A(KEYINPUT97), .ZN(n656) );
  INV_X1 U567 ( .A(KEYINPUT101), .ZN(n701) );
  XNOR2_X1 U568 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U569 ( .A1(n714), .A2(n603), .ZN(n666) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n590) );
  INV_X1 U571 ( .A(KEYINPUT9), .ZN(n568) );
  AND2_X2 U572 ( .A1(n524), .A2(G2104), .ZN(n895) );
  INV_X1 U573 ( .A(KEYINPUT23), .ZN(n525) );
  XNOR2_X1 U574 ( .A(KEYINPUT66), .B(n544), .ZN(n806) );
  XNOR2_X1 U575 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U576 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n524), .ZN(n890) );
  NAND2_X1 U579 ( .A1(n890), .A2(G125), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G101), .A2(n895), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n534) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n530), .B(n529), .ZN(n715) );
  NAND2_X1 U585 ( .A1(G137), .A2(n715), .ZN(n532) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U587 ( .A1(G113), .A2(n891), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n802) );
  NAND2_X1 U590 ( .A1(G89), .A2(n802), .ZN(n535) );
  XOR2_X1 U591 ( .A(KEYINPUT4), .B(n535), .Z(n536) );
  XNOR2_X1 U592 ( .A(n536), .B(KEYINPUT75), .ZN(n539) );
  INV_X1 U593 ( .A(G651), .ZN(n541) );
  OR2_X1 U594 ( .A1(n541), .A2(n590), .ZN(n537) );
  XOR2_X2 U595 ( .A(KEYINPUT68), .B(n537), .Z(n805) );
  NAND2_X1 U596 ( .A1(G76), .A2(n805), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n540), .B(KEYINPUT5), .ZN(n549) );
  NOR2_X1 U599 ( .A1(G543), .A2(n541), .ZN(n543) );
  XNOR2_X1 U600 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n543), .B(n542), .ZN(n801) );
  NAND2_X1 U602 ( .A1(G63), .A2(n801), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n590), .A2(G651), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G51), .A2(n806), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U606 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G138), .A2(n715), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G102), .A2(n895), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G126), .A2(n890), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G114), .A2(n891), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U615 ( .A1(G65), .A2(n801), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G91), .A2(n802), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G78), .A2(n805), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G53), .A2(n806), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G299) );
  NAND2_X1 U622 ( .A1(G64), .A2(n801), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G52), .A2(n806), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G77), .A2(n805), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT71), .B(n565), .Z(n567) );
  NAND2_X1 U627 ( .A1(n802), .A2(G90), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n569) );
  NOR2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U630 ( .A(KEYINPUT72), .B(n572), .ZN(G171) );
  NAND2_X1 U631 ( .A1(G88), .A2(n802), .ZN(n573) );
  XNOR2_X1 U632 ( .A(n573), .B(KEYINPUT82), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n805), .A2(G75), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT83), .B(n574), .Z(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G62), .A2(n801), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G50), .A2(n806), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U639 ( .A1(n580), .A2(n579), .ZN(G166) );
  XNOR2_X1 U640 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G61), .A2(n801), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G86), .A2(n802), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n805), .A2(G73), .ZN(n583) );
  XNOR2_X1 U646 ( .A(n583), .B(KEYINPUT81), .ZN(n584) );
  XNOR2_X1 U647 ( .A(n584), .B(KEYINPUT2), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U649 ( .A1(G48), .A2(n806), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G74), .A2(G651), .ZN(n589) );
  XNOR2_X1 U652 ( .A(n589), .B(KEYINPUT80), .ZN(n595) );
  NAND2_X1 U653 ( .A1(n590), .A2(G87), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G49), .A2(n806), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U656 ( .A1(n801), .A2(n593), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(G288) );
  NAND2_X1 U658 ( .A1(n802), .A2(G85), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n801), .A2(G60), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U661 ( .A1(G72), .A2(n805), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G47), .A2(n806), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U664 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U665 ( .A(KEYINPUT70), .B(n602), .Z(G290) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n714) );
  NAND2_X1 U667 ( .A1(G160), .A2(G40), .ZN(n713) );
  INV_X1 U668 ( .A(n713), .ZN(n603) );
  NOR2_X1 U669 ( .A1(G2084), .A2(n666), .ZN(n651) );
  NAND2_X1 U670 ( .A1(n651), .A2(G8), .ZN(n665) );
  NAND2_X1 U671 ( .A1(G8), .A2(n666), .ZN(n706) );
  NOR2_X1 U672 ( .A1(G1966), .A2(n706), .ZN(n663) );
  INV_X1 U673 ( .A(KEYINPUT93), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(n646), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n607), .A2(G2072), .ZN(n605) );
  INV_X1 U676 ( .A(n607), .ZN(n645) );
  NAND2_X1 U677 ( .A1(G1956), .A2(n645), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n523), .A2(n606), .ZN(n640) );
  NOR2_X1 U679 ( .A1(G299), .A2(n640), .ZN(n619) );
  NAND2_X1 U680 ( .A1(G2067), .A2(n607), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G1348), .A2(n666), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT94), .ZN(n620) );
  NAND2_X1 U684 ( .A1(G79), .A2(n805), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G54), .A2(n806), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G66), .A2(n801), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G92), .A2(n802), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT15), .ZN(n990) );
  NOR2_X1 U692 ( .A1(n620), .A2(n990), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n638) );
  NAND2_X1 U694 ( .A1(n990), .A2(n620), .ZN(n636) );
  NAND2_X1 U695 ( .A1(G56), .A2(n801), .ZN(n621) );
  XOR2_X1 U696 ( .A(KEYINPUT14), .B(n621), .Z(n627) );
  NAND2_X1 U697 ( .A1(n802), .A2(G81), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n622), .B(KEYINPUT12), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G68), .A2(n805), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U701 ( .A(KEYINPUT13), .B(n625), .Z(n626) );
  NOR2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G43), .A2(n806), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n1002) );
  INV_X1 U705 ( .A(G1996), .ZN(n963) );
  NOR2_X1 U706 ( .A1(n666), .A2(n963), .ZN(n631) );
  XNOR2_X1 U707 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n631), .B(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n666), .A2(G1341), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n1002), .A2(n634), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  AND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n639), .B(KEYINPUT95), .ZN(n643) );
  NAND2_X1 U715 ( .A1(G299), .A2(n640), .ZN(n641) );
  XNOR2_X1 U716 ( .A(KEYINPUT28), .B(n641), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(KEYINPUT29), .ZN(n675) );
  INV_X1 U719 ( .A(G171), .ZN(n650) );
  XOR2_X1 U720 ( .A(KEYINPUT25), .B(G2078), .Z(n964) );
  NOR2_X1 U721 ( .A1(n964), .A2(n645), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n646), .A2(G1961), .ZN(n647) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n673) );
  NOR2_X1 U725 ( .A1(n675), .A2(n673), .ZN(n661) );
  AND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n663), .A2(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G8), .A2(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U731 ( .A1(G168), .A2(n655), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(KEYINPUT31), .ZN(n677) );
  NOR2_X1 U735 ( .A1(n661), .A2(n677), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n685) );
  INV_X1 U738 ( .A(G8), .ZN(n671) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n706), .ZN(n668) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n666), .ZN(n667) );
  NOR2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(G303), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n676) );
  OR2_X1 U744 ( .A1(n676), .A2(G286), .ZN(n679) );
  INV_X1 U745 ( .A(n679), .ZN(n672) );
  NOR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n699) );
  INV_X1 U749 ( .A(n699), .ZN(n689) );
  NOR2_X1 U750 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U751 ( .A1(G8), .A2(n686), .ZN(n687) );
  XOR2_X1 U752 ( .A(KEYINPUT102), .B(n687), .Z(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(KEYINPUT103), .B(n690), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n691), .A2(n706), .ZN(n759) );
  NOR2_X1 U756 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XOR2_X1 U757 ( .A(n692), .B(KEYINPUT24), .Z(n693) );
  NOR2_X1 U758 ( .A1(n706), .A2(n693), .ZN(n712) );
  NOR2_X1 U759 ( .A1(G288), .A2(G1976), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(KEYINPUT99), .ZN(n993) );
  INV_X1 U761 ( .A(n993), .ZN(n696) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT100), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NAND2_X1 U767 ( .A1(n700), .A2(n994), .ZN(n702) );
  NOR2_X1 U768 ( .A1(n703), .A2(n706), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT64), .ZN(n705) );
  NOR2_X1 U770 ( .A1(KEYINPUT33), .A2(n705), .ZN(n710) );
  NOR2_X1 U771 ( .A1(n706), .A2(n993), .ZN(n707) );
  NAND2_X1 U772 ( .A1(KEYINPUT33), .A2(n707), .ZN(n708) );
  XOR2_X1 U773 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U774 ( .A1(n708), .A2(n983), .ZN(n709) );
  NOR2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n759), .A2(n761), .ZN(n747) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n765) );
  XNOR2_X1 U778 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NAND2_X1 U779 ( .A1(G140), .A2(n716), .ZN(n718) );
  NAND2_X1 U780 ( .A1(G104), .A2(n895), .ZN(n717) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n720) );
  XOR2_X1 U782 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n719) );
  XNOR2_X1 U783 ( .A(n720), .B(n719), .ZN(n726) );
  NAND2_X1 U784 ( .A1(n891), .A2(G116), .ZN(n721) );
  XNOR2_X1 U785 ( .A(n721), .B(KEYINPUT92), .ZN(n723) );
  NAND2_X1 U786 ( .A1(G128), .A2(n890), .ZN(n722) );
  NAND2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U788 ( .A(KEYINPUT35), .B(n724), .Z(n725) );
  NOR2_X1 U789 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U790 ( .A(KEYINPUT36), .B(n727), .ZN(n907) );
  NOR2_X1 U791 ( .A1(n753), .A2(n907), .ZN(n951) );
  NAND2_X1 U792 ( .A1(n765), .A2(n951), .ZN(n764) );
  XNOR2_X1 U793 ( .A(G1986), .B(G290), .ZN(n989) );
  AND2_X1 U794 ( .A1(n989), .A2(n765), .ZN(n744) );
  NAND2_X1 U795 ( .A1(G141), .A2(n716), .ZN(n729) );
  NAND2_X1 U796 ( .A1(G129), .A2(n890), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U798 ( .A1(n895), .A2(G105), .ZN(n730) );
  XOR2_X1 U799 ( .A(KEYINPUT38), .B(n730), .Z(n731) );
  NOR2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U801 ( .A1(n891), .A2(G117), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n903) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n903), .ZN(n742) );
  NAND2_X1 U804 ( .A1(G131), .A2(n716), .ZN(n736) );
  NAND2_X1 U805 ( .A1(G119), .A2(n890), .ZN(n735) );
  NAND2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n740) );
  NAND2_X1 U807 ( .A1(G95), .A2(n895), .ZN(n738) );
  NAND2_X1 U808 ( .A1(G107), .A2(n891), .ZN(n737) );
  NAND2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n887) );
  NAND2_X1 U811 ( .A1(G1991), .A2(n887), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n947) );
  NAND2_X1 U813 ( .A1(n765), .A2(n947), .ZN(n748) );
  NAND2_X1 U814 ( .A1(KEYINPUT90), .A2(n748), .ZN(n743) );
  NOR2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U816 ( .A1(n764), .A2(n745), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n747), .A2(n746), .ZN(n774) );
  INV_X1 U818 ( .A(n765), .ZN(n758) );
  INV_X1 U819 ( .A(n764), .ZN(n756) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n903), .ZN(n938) );
  INV_X1 U821 ( .A(n748), .ZN(n763) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n749) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n887), .ZN(n944) );
  NOR2_X1 U824 ( .A1(n749), .A2(n944), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n763), .A2(n750), .ZN(n751) );
  NOR2_X1 U826 ( .A1(n938), .A2(n751), .ZN(n752) );
  XOR2_X1 U827 ( .A(KEYINPUT39), .B(n752), .Z(n754) );
  NAND2_X1 U828 ( .A1(n753), .A2(n907), .ZN(n956) );
  AND2_X1 U829 ( .A1(n754), .A2(n956), .ZN(n755) );
  OR2_X1 U830 ( .A1(n756), .A2(n755), .ZN(n757) );
  OR2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n762) );
  AND2_X1 U832 ( .A1(n759), .A2(n762), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n772) );
  INV_X1 U834 ( .A(n762), .ZN(n770) );
  NOR2_X1 U835 ( .A1(KEYINPUT90), .A2(n763), .ZN(n768) );
  AND2_X1 U836 ( .A1(n989), .A2(n764), .ZN(n766) );
  AND2_X1 U837 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U838 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U839 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U840 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U841 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U842 ( .A(n775), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  INV_X1 U846 ( .A(G120), .ZN(G236) );
  INV_X1 U847 ( .A(G69), .ZN(G235) );
  INV_X1 U848 ( .A(G108), .ZN(G238) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U850 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U851 ( .A(G223), .ZN(n838) );
  NAND2_X1 U852 ( .A1(n838), .A2(G567), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n777), .B(KEYINPUT73), .ZN(n778) );
  XNOR2_X1 U854 ( .A(KEYINPUT11), .B(n778), .ZN(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n845) );
  OR2_X1 U856 ( .A1(n1002), .A2(n845), .ZN(G153) );
  XNOR2_X1 U857 ( .A(n650), .B(KEYINPUT74), .ZN(G301) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n780) );
  INV_X1 U859 ( .A(G868), .ZN(n819) );
  NAND2_X1 U860 ( .A1(n990), .A2(n819), .ZN(n779) );
  NAND2_X1 U861 ( .A1(n780), .A2(n779), .ZN(G284) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n782) );
  NOR2_X1 U863 ( .A1(G286), .A2(n819), .ZN(n781) );
  NOR2_X1 U864 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U865 ( .A1(n845), .A2(G559), .ZN(n783) );
  INV_X1 U866 ( .A(n990), .ZN(n799) );
  NAND2_X1 U867 ( .A1(n783), .A2(n799), .ZN(n784) );
  XNOR2_X1 U868 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U869 ( .A1(G868), .A2(n1002), .ZN(n787) );
  NAND2_X1 U870 ( .A1(G868), .A2(n799), .ZN(n785) );
  NOR2_X1 U871 ( .A1(G559), .A2(n785), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(G282) );
  XOR2_X1 U873 ( .A(G2100), .B(KEYINPUT78), .Z(n798) );
  NAND2_X1 U874 ( .A1(n890), .A2(G123), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n788), .B(KEYINPUT18), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G135), .A2(n716), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U878 ( .A(KEYINPUT76), .B(n791), .Z(n793) );
  NAND2_X1 U879 ( .A1(n891), .A2(G111), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G99), .A2(n895), .ZN(n794) );
  XNOR2_X1 U882 ( .A(KEYINPUT77), .B(n794), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n943) );
  XNOR2_X1 U884 ( .A(G2096), .B(n943), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G559), .A2(n799), .ZN(n800) );
  XOR2_X1 U887 ( .A(n1002), .B(n800), .Z(n844) );
  NAND2_X1 U888 ( .A1(G67), .A2(n801), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n810) );
  NAND2_X1 U891 ( .A1(G80), .A2(n805), .ZN(n808) );
  NAND2_X1 U892 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U895 ( .A(KEYINPUT79), .B(n811), .ZN(n846) );
  XOR2_X1 U896 ( .A(G299), .B(n846), .Z(n813) );
  XNOR2_X1 U897 ( .A(G290), .B(G166), .ZN(n812) );
  XNOR2_X1 U898 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U899 ( .A(n814), .B(G305), .ZN(n817) );
  XNOR2_X1 U900 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n815), .B(G288), .ZN(n816) );
  XNOR2_X1 U902 ( .A(n817), .B(n816), .ZN(n911) );
  XNOR2_X1 U903 ( .A(n844), .B(n911), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n818), .A2(G868), .ZN(n821) );
  NAND2_X1 U905 ( .A1(n819), .A2(n846), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n821), .A2(n820), .ZN(G295) );
  XOR2_X1 U907 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n825) );
  NAND2_X1 U908 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U910 ( .A1(n823), .A2(G2090), .ZN(n824) );
  XNOR2_X1 U911 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U912 ( .A(KEYINPUT86), .B(n826), .ZN(n827) );
  NAND2_X1 U913 ( .A1(n827), .A2(G2072), .ZN(n828) );
  XOR2_X1 U914 ( .A(KEYINPUT87), .B(n828), .Z(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G235), .A2(G236), .ZN(n829) );
  XOR2_X1 U917 ( .A(KEYINPUT88), .B(n829), .Z(n830) );
  NOR2_X1 U918 ( .A1(G238), .A2(n830), .ZN(n831) );
  NAND2_X1 U919 ( .A1(G57), .A2(n831), .ZN(n842) );
  NAND2_X1 U920 ( .A1(n842), .A2(G567), .ZN(n836) );
  NOR2_X1 U921 ( .A1(G220), .A2(G219), .ZN(n832) );
  XOR2_X1 U922 ( .A(KEYINPUT22), .B(n832), .Z(n833) );
  NOR2_X1 U923 ( .A1(G218), .A2(n833), .ZN(n834) );
  NAND2_X1 U924 ( .A1(G96), .A2(n834), .ZN(n843) );
  NAND2_X1 U925 ( .A1(n843), .A2(G2106), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n836), .A2(n835), .ZN(n848) );
  NAND2_X1 U927 ( .A1(G483), .A2(G661), .ZN(n837) );
  NOR2_X1 U928 ( .A1(n848), .A2(n837), .ZN(n841) );
  NAND2_X1 U929 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U932 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n841), .A2(n840), .ZN(G188) );
  NOR2_X1 U935 ( .A1(n843), .A2(n842), .ZN(G325) );
  XOR2_X1 U936 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(n847) );
  XNOR2_X1 U940 ( .A(n847), .B(n846), .ZN(G145) );
  INV_X1 U941 ( .A(n848), .ZN(G319) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G1991), .Z(n850) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1981), .ZN(n849) );
  XNOR2_X1 U944 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U945 ( .A(n851), .B(KEYINPUT109), .Z(n853) );
  XNOR2_X1 U946 ( .A(G1971), .B(G1956), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U948 ( .A(G1976), .B(G1966), .Z(n855) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1961), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U951 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U952 ( .A(KEYINPUT108), .B(G2474), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n859), .B(n858), .ZN(G229) );
  XOR2_X1 U954 ( .A(KEYINPUT107), .B(G2084), .Z(n861) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2090), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U957 ( .A(n862), .B(G2096), .Z(n864) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2072), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U960 ( .A(G2100), .B(G2678), .Z(n866) );
  XNOR2_X1 U961 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U963 ( .A(n868), .B(n867), .Z(G227) );
  NAND2_X1 U964 ( .A1(G124), .A2(n890), .ZN(n869) );
  XNOR2_X1 U965 ( .A(n869), .B(KEYINPUT44), .ZN(n870) );
  XNOR2_X1 U966 ( .A(n870), .B(KEYINPUT110), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G112), .A2(n891), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G136), .A2(n716), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G100), .A2(n895), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U972 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G139), .A2(n716), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G103), .A2(n895), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U976 ( .A1(G127), .A2(n890), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G115), .A2(n891), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n933) );
  XOR2_X1 U981 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n933), .B(n886), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n887), .B(n943), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n902) );
  NAND2_X1 U987 ( .A1(G130), .A2(n890), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U990 ( .A1(n716), .A2(G142), .ZN(n894) );
  XOR2_X1 U991 ( .A(KEYINPUT111), .B(n894), .Z(n897) );
  NAND2_X1 U992 ( .A1(n895), .A2(G106), .ZN(n896) );
  NAND2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(n902), .B(n901), .Z(n909) );
  XNOR2_X1 U997 ( .A(n903), .B(G162), .ZN(n905) );
  XNOR2_X1 U998 ( .A(G164), .B(G160), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1000 ( .A(n907), .B(n906), .Z(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n911), .B(n1002), .ZN(n912) );
  XNOR2_X1 U1004 ( .A(n912), .B(n990), .ZN(n914) );
  XOR2_X1 U1005 ( .A(G171), .B(G286), .Z(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n915), .ZN(G397) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2443), .ZN(n925) );
  XOR2_X1 U1009 ( .A(G2446), .B(G2430), .Z(n917) );
  XNOR2_X1 U1010 ( .A(KEYINPUT105), .B(G2438), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n921) );
  XOR2_X1 U1012 ( .A(G2435), .B(G2454), .Z(n919) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1015 ( .A(n921), .B(n920), .Z(n923) );
  XNOR2_X1 U1016 ( .A(KEYINPUT104), .B(G2427), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1019 ( .A1(n926), .A2(G14), .ZN(n932) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n932), .ZN(n929) );
  NOR2_X1 U1021 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G57), .ZN(G237) );
  INV_X1 U1028 ( .A(n932), .ZN(G401) );
  XNOR2_X1 U1029 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1043) );
  INV_X1 U1030 ( .A(KEYINPUT55), .ZN(n960) );
  XOR2_X1 U1031 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(KEYINPUT50), .B(n936), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  XNOR2_X1 U1038 ( .A(KEYINPUT116), .B(n940), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n954) );
  XNOR2_X1 U1040 ( .A(G160), .B(G2084), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1042 ( .A(KEYINPUT114), .B(n945), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT115), .B(n952), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(n957), .B(KEYINPUT117), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n958), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1052 ( .A1(n961), .A2(G29), .ZN(n1041) );
  XNOR2_X1 U1053 ( .A(G2084), .B(G34), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n962), .B(KEYINPUT54), .ZN(n980) );
  XOR2_X1 U1055 ( .A(G2090), .B(G35), .Z(n978) );
  XNOR2_X1 U1056 ( .A(G32), .B(n963), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G27), .B(n964), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(G33), .B(G2072), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1063 ( .A(KEYINPUT118), .B(n971), .Z(n973) );
  XNOR2_X1 U1064 ( .A(G1991), .B(G25), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n974), .A2(G28), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT53), .B(n975), .Z(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT119), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1071 ( .A(KEYINPUT55), .B(n981), .Z(n982) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n982), .ZN(n1037) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1074 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n985), .B(KEYINPUT57), .ZN(n1006) );
  XNOR2_X1 U1077 ( .A(G303), .B(G1971), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(n650), .B(G1961), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n1000) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G299), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1082 ( .A(G1348), .B(n990), .Z(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT120), .B(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1086 ( .A(KEYINPUT121), .B(n996), .Z(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(KEYINPUT122), .B(n1001), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1035) );
  INV_X1 U1094 ( .A(G16), .ZN(n1033) );
  XOR2_X1 U1095 ( .A(G1976), .B(G23), .Z(n1010) );
  XOR2_X1 U1096 ( .A(G1971), .B(G22), .Z(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G24), .B(G1986), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1013), .Z(n1030) );
  XOR2_X1 U1101 ( .A(G1961), .B(G5), .Z(n1025) );
  XNOR2_X1 U1102 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(n1014), .B(G4), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G1348), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G1341), .B(G19), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(G1956), .B(G20), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(KEYINPUT124), .B(n1022), .Z(n1023) );
  XNOR2_X1 U1112 ( .A(n1023), .B(KEYINPUT60), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(G21), .B(G1966), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT125), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1122 ( .A1(G11), .A2(n1038), .ZN(n1039) );
  XOR2_X1 U1123 ( .A(KEYINPUT126), .B(n1039), .Z(n1040) );
  NAND2_X1 U1124 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1125 ( .A(n1043), .B(n1042), .ZN(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

