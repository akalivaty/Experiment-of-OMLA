//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT0), .A3(G128), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G128), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n187), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT11), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT64), .A2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n195), .A2(new_n196), .A3(new_n200), .A4(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT11), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n196), .B1(new_n203), .B2(new_n194), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n192), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(G131), .ZN(new_n207));
  AOI211_X1 g021(.A(new_n207), .B(new_n204), .C1(new_n199), .C2(new_n201), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n191), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT70), .A2(G116), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT70), .A2(G116), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n216), .B2(G119), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n211), .B1(new_n217), .B2(KEYINPUT69), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n214), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n219), .B(new_n210), .C1(new_n221), .C2(new_n213), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n207), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT64), .A2(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT64), .A2(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n200), .B1(new_n228), .B2(new_n196), .ZN(new_n229));
  INV_X1    g043(.A(new_n201), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n225), .B(new_n205), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G128), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n233), .B(new_n235), .C1(KEYINPUT1), .C2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n228), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G131), .C1(new_n242), .C2(new_n194), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n209), .A2(new_n224), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n224), .B1(new_n209), .B2(new_n245), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT28), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT73), .ZN(new_n250));
  INV_X1    g064(.A(G237), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT71), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G237), .ZN(new_n254));
  AOI21_X1  g068(.A(G953), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n250), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n257), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n209), .A2(new_n245), .A3(new_n224), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n248), .A2(KEYINPUT29), .A3(new_n260), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n260), .A2(new_n263), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n205), .B1(new_n229), .B2(new_n230), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  AOI211_X1 g086(.A(KEYINPUT67), .B(new_n190), .C1(new_n272), .C2(new_n231), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n204), .B1(new_n199), .B2(new_n201), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n231), .B1(new_n192), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n276), .B2(new_n191), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n245), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n246), .B1(new_n278), .B2(new_n223), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n270), .B1(new_n279), .B2(new_n262), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT75), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n270), .B(new_n283), .C1(new_n279), .C2(new_n262), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n231), .A2(new_n241), .A3(new_n244), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n276), .B2(new_n191), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT30), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n223), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n274), .A3(new_n191), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT30), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT68), .B1(new_n278), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n290), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n260), .B1(new_n298), .B2(new_n261), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n269), .B1(new_n285), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G472), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  INV_X1    g116(.A(new_n260), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(new_n246), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n263), .B1(new_n279), .B2(new_n262), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n294), .B1(new_n293), .B2(KEYINPUT30), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n278), .A2(KEYINPUT68), .A3(new_n296), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n289), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n304), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT74), .B1(new_n313), .B2(new_n302), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n315), .B(KEYINPUT31), .C1(new_n311), .C2(new_n312), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n308), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G472), .A2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n301), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n313), .A2(new_n302), .B1(new_n303), .B2(new_n306), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n298), .A2(new_n304), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n315), .B1(new_n325), .B2(KEYINPUT31), .ZN(new_n326));
  INV_X1    g140(.A(new_n316), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT32), .B1(new_n328), .B2(new_n318), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT77), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n328), .A2(new_n321), .B1(new_n300), .B2(G472), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n320), .B1(new_n317), .B2(new_n319), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT16), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G125), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT80), .A4(G125), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n342));
  AND3_X1   g156(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n343));
  AOI21_X1  g157(.A(G140), .B1(KEYINPUT79), .B2(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT16), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n341), .A2(new_n342), .A3(G146), .A4(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(G146), .A3(new_n339), .A4(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT81), .ZN(new_n348));
  INV_X1    g162(.A(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n339), .A2(new_n340), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n232), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n220), .B2(G128), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n354), .B(new_n355), .C1(G119), .C2(new_n239), .ZN(new_n356));
  XNOR2_X1  g170(.A(G119), .B(G128), .ZN(new_n357));
  XOR2_X1   g171(.A(KEYINPUT24), .B(G110), .Z(new_n358));
  AOI22_X1  g172(.A1(new_n356), .A2(G110), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G125), .B(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n232), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT82), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(new_n232), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI22_X1  g180(.A1(new_n356), .A2(G110), .B1(new_n357), .B2(new_n358), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n347), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(G221), .A3(G234), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT83), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G137), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n360), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n360), .B2(new_n368), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n266), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g191(.A1(G217), .A2(G902), .ZN(new_n378));
  INV_X1    g192(.A(G217), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(G234), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT78), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT25), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n266), .C1(new_n374), .C2(new_n375), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n374), .A2(new_n375), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n381), .A2(G902), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G469), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G104), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G107), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n396), .B2(new_n394), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT86), .B(G101), .Z(new_n398));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(G104), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(KEYINPUT3), .C1(new_n393), .C2(G107), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n397), .B(new_n398), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n241), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT10), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n390), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n395), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n408), .A2(KEYINPUT87), .A3(KEYINPUT10), .A4(new_n241), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n276), .ZN(new_n411));
  INV_X1    g225(.A(G101), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n393), .A2(G107), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT85), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n416), .B2(new_n402), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n404), .B(KEYINPUT4), .C1(new_n412), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n402), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n412), .B1(new_n419), .B2(new_n397), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n190), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n418), .A2(new_n422), .B1(new_n405), .B2(new_n406), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(new_n411), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  INV_X1    g239(.A(G227), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n425), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n404), .A2(new_n395), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n238), .A2(new_n240), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n405), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT12), .A3(new_n276), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT12), .B1(new_n433), .B2(new_n276), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n424), .B(new_n429), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n410), .A2(new_n423), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n276), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n429), .B1(new_n440), .B2(new_n424), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n389), .B(new_n266), .C1(new_n438), .C2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n389), .A2(new_n266), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n435), .A2(new_n436), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n410), .A2(new_n411), .A3(new_n423), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n428), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n424), .A2(new_n448), .A3(new_n429), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n440), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n424), .B2(new_n429), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n447), .B(G469), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n444), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT9), .B(G234), .ZN(new_n455));
  OAI21_X1  g269(.A(G221), .B1(new_n455), .B2(G902), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT84), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n454), .B1(new_n453), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G214), .B1(G237), .B2(G902), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT90), .ZN(new_n463));
  INV_X1    g277(.A(G125), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n238), .A2(new_n464), .A3(new_n240), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n190), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n369), .A2(G224), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(KEYINPUT7), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT94), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(KEYINPUT7), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n465), .B(new_n470), .C1(new_n190), .C2(new_n464), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT93), .Z(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT8), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g289(.A(new_n213), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(G113), .C1(KEYINPUT5), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n217), .A2(new_n211), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n477), .A2(new_n408), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n408), .B1(new_n478), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(new_n472), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n420), .A2(new_n421), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n418), .A2(new_n223), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n222), .A2(new_n218), .B1(new_n420), .B2(new_n421), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n418), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n477), .A2(new_n408), .A3(new_n478), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(new_n473), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n266), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  AND2_X1   g308(.A1(KEYINPUT92), .A2(KEYINPUT6), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n473), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(new_n489), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n487), .B1(new_n486), .B2(new_n418), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n497), .B(new_n495), .C1(new_n498), .C2(new_n499), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n466), .B(new_n467), .Z(new_n504));
  OAI211_X1 g318(.A(new_n493), .B(new_n494), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n494), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n504), .B1(new_n501), .B2(new_n502), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n492), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n463), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n369), .A2(G952), .ZN(new_n510));
  INV_X1    g324(.A(G234), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n251), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n266), .B(new_n369), .C1(G234), .C2(G237), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G113), .B(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n393), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT95), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n252), .A2(new_n254), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(G214), .A3(new_n369), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n234), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT18), .A3(G131), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n343), .A2(new_n344), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G146), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n366), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT18), .A2(G131), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n207), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n225), .A3(new_n524), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n525), .A2(KEYINPUT17), .A3(new_n207), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n538), .A2(new_n348), .A3(new_n351), .A4(new_n346), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n520), .B(new_n532), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n266), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n534), .B(new_n225), .C1(new_n523), .C2(new_n524), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n352), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n520), .B1(new_n544), .B2(new_n532), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT96), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n532), .B1(new_n537), .B2(new_n539), .ZN(new_n547));
  INV_X1    g361(.A(new_n520), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n266), .A4(new_n540), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(G475), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n519), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n533), .A2(new_n535), .ZN(new_n554));
  MUX2_X1   g368(.A(new_n361), .B(new_n527), .S(KEYINPUT19), .Z(new_n555));
  OAI21_X1  g369(.A(new_n347), .B1(new_n555), .B2(G146), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n553), .B(new_n532), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n529), .A2(new_n531), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n543), .A2(new_n536), .B1(new_n559), .B2(new_n526), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n557), .B(new_n558), .C1(new_n560), .C2(new_n553), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT20), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n547), .A2(new_n519), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n557), .A4(new_n558), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n552), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n455), .A2(new_n379), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT13), .B1(new_n239), .B2(G143), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n242), .ZN(new_n571));
  XNOR2_X1  g385(.A(G128), .B(G143), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(KEYINPUT98), .ZN(new_n574));
  OR2_X1    g388(.A1(KEYINPUT70), .A2(G116), .ZN(new_n575));
  NAND2_X1  g389(.A1(KEYINPUT70), .A2(G116), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(G122), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n212), .A2(G122), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n578), .B1(new_n577), .B2(new_n580), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n582), .A2(new_n583), .A3(new_n391), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT97), .ZN(new_n586));
  AOI21_X1  g400(.A(G107), .B1(new_n586), .B2(new_n581), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n574), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n391), .B1(new_n582), .B2(new_n583), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n581), .A3(G107), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT98), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n573), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n572), .B(new_n242), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n585), .A2(KEYINPUT14), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT14), .ZN(new_n595));
  OAI21_X1  g409(.A(G107), .B1(new_n577), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n593), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n587), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n569), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n573), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n589), .A2(KEYINPUT98), .A3(new_n590), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT98), .B1(new_n589), .B2(new_n590), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n598), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n568), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n266), .ZN(new_n607));
  INV_X1    g421(.A(G478), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(KEYINPUT15), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(new_n266), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n567), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n509), .A2(new_n517), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n461), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n330), .A2(new_n334), .A3(new_n388), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(new_n398), .Z(G3));
  NAND2_X1  g432(.A1(new_n328), .A2(new_n266), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n328), .A2(new_n318), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n388), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n461), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n509), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n607), .A2(G478), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n608), .A2(new_n266), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(G478), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n567), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n625), .A2(new_n516), .A3(new_n626), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT100), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  NAND2_X1  g453(.A1(new_n505), .A2(new_n508), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n611), .B1(new_n606), .B2(new_n266), .ZN(new_n641));
  AOI211_X1 g455(.A(G902), .B(new_n609), .C1(new_n599), .C2(new_n605), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n567), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n463), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n640), .A2(new_n644), .A3(new_n517), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT101), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n622), .A2(new_n624), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NAND2_X1  g464(.A1(new_n360), .A2(new_n368), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n373), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n386), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n384), .A2(KEYINPUT102), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT102), .B1(new_n384), .B2(new_n654), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n622), .A2(new_n616), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n509), .A2(new_n658), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n461), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n644), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n514), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n512), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n330), .A2(new_n334), .A3(new_n663), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XNOR2_X1  g485(.A(new_n640), .B(KEYINPUT38), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n567), .A2(new_n613), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n463), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n667), .B(KEYINPUT39), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n459), .B2(new_n460), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n672), .B(new_n674), .C1(new_n676), .C2(KEYINPUT40), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(KEYINPUT40), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n384), .A2(new_n654), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n303), .B1(new_n246), .B2(new_n247), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n325), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n266), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n328), .A2(new_n321), .B1(G472), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT103), .B1(new_n332), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n332), .A2(new_n684), .A3(KEYINPUT103), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n678), .B(new_n680), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NAND3_X1  g502(.A1(new_n633), .A2(new_n567), .A3(new_n667), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n461), .A2(new_n662), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n330), .A2(new_n334), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n330), .A2(new_n690), .A3(KEYINPUT104), .A4(new_n334), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NOR2_X1   g510(.A1(new_n389), .A2(KEYINPUT105), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n411), .B1(new_n410), .B2(new_n423), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n428), .B1(new_n446), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n437), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n701), .B2(new_n266), .ZN(new_n702));
  AOI211_X1 g516(.A(G902), .B(new_n697), .C1(new_n700), .C2(new_n437), .ZN(new_n703));
  INV_X1    g517(.A(new_n456), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n623), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n634), .A2(new_n626), .A3(new_n516), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n330), .A2(new_n334), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n330), .A2(new_n647), .A3(new_n334), .A4(new_n707), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NOR2_X1   g527(.A1(new_n626), .A2(new_n706), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n658), .A2(new_n517), .A3(new_n614), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n330), .A2(new_n334), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  XNOR2_X1  g531(.A(KEYINPUT106), .B(G472), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n317), .B2(G902), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n567), .A2(new_n517), .A3(new_n613), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n509), .A2(new_n720), .A3(new_n705), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n260), .B1(new_n248), .B2(new_n263), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n313), .B2(new_n302), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n325), .A2(KEYINPUT31), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n319), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n719), .A2(new_n721), .A3(new_n388), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n725), .B1(new_n619), .B2(new_n718), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(KEYINPUT107), .A3(new_n388), .A4(new_n721), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  INV_X1    g547(.A(new_n689), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n679), .A3(new_n734), .A4(new_n714), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(new_n447), .ZN(new_n737));
  OR3_X1    g551(.A1(new_n450), .A2(KEYINPUT108), .A3(new_n451), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT108), .B1(new_n450), .B2(new_n451), .ZN(new_n739));
  AOI211_X1 g553(.A(new_n389), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n442), .A2(new_n444), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n456), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n505), .A2(new_n645), .A3(new_n508), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n742), .A2(new_n689), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n623), .B1(new_n331), .B2(new_n332), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n330), .A2(new_n334), .A3(new_n388), .A4(new_n744), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(KEYINPUT109), .A3(new_n746), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT109), .B1(new_n750), .B2(new_n746), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  AND3_X1   g569(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n742), .A2(new_n743), .A3(new_n623), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n669), .A4(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n330), .A2(new_n334), .A3(new_n669), .A4(new_n760), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  INV_X1    g579(.A(new_n622), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n633), .A2(new_n552), .A3(new_n566), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT43), .Z(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n679), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n743), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n389), .B(new_n774), .C1(new_n775), .C2(KEYINPUT45), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n443), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n442), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n456), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n675), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n771), .B(new_n782), .C1(new_n770), .C2(new_n769), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  XOR2_X1   g598(.A(new_n780), .B(KEYINPUT47), .Z(new_n785));
  NOR4_X1   g599(.A1(new_n758), .A2(new_n388), .A3(new_n689), .A4(new_n743), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n388), .A2(new_n458), .A3(new_n645), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n767), .B1(KEYINPUT111), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(KEYINPUT111), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n702), .A2(new_n703), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT49), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT49), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n791), .A2(new_n792), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n672), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n686), .A2(new_n685), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n617), .A2(new_n732), .A3(new_n709), .A4(new_n712), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n744), .A2(new_n679), .A3(new_n730), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n658), .A2(new_n614), .A3(new_n667), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n461), .A2(new_n743), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n330), .A2(new_n334), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT112), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n330), .A2(new_n804), .A3(new_n807), .A4(new_n334), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n802), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n626), .A2(new_n516), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n634), .A2(new_n664), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n622), .A2(new_n810), .A3(new_n624), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n716), .A3(new_n659), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n801), .A2(new_n764), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n750), .A2(new_n746), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n818), .A2(new_n751), .B1(new_n748), .B2(new_n747), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n764), .A2(new_n809), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n732), .A2(new_n712), .A3(new_n617), .A4(new_n709), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n813), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n754), .A4(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n670), .A2(new_n735), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n742), .A2(new_n626), .A3(new_n668), .A4(new_n673), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n680), .B(new_n827), .C1(new_n686), .C2(new_n685), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n695), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n695), .A2(new_n826), .A3(KEYINPUT52), .A4(new_n828), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n834), .A3(new_n830), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n820), .A2(new_n825), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT115), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n821), .A2(new_n754), .A3(new_n824), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n831), .A2(new_n832), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n832), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n839), .A2(new_n841), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n768), .A2(new_n513), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n730), .A2(new_n388), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n672), .A2(new_n706), .A3(new_n645), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT50), .Z(new_n855));
  NOR2_X1   g669(.A1(new_n706), .A2(new_n743), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n799), .A2(new_n388), .A3(new_n513), .A4(new_n856), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n857), .A2(new_n567), .A3(new_n633), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n768), .A2(new_n513), .A3(new_n856), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n679), .A3(new_n730), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n855), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n850), .A2(new_n851), .A3(new_n743), .ZN(new_n863));
  INV_X1    g677(.A(new_n785), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n793), .A2(new_n457), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT117), .Z(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT51), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n862), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n860), .A2(new_n748), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT48), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n852), .A2(new_n714), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n875), .B(new_n510), .C1(new_n634), .C2(new_n857), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n869), .A2(new_n872), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n845), .B2(new_n846), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n815), .A2(new_n819), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n833), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n849), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n789), .B(new_n800), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n878), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n848), .B2(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n889), .B2(new_n877), .ZN(new_n890));
  INV_X1    g704(.A(new_n800), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT119), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n882), .A2(new_n266), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G210), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n503), .B(new_n504), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n369), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  NAND2_X1  g716(.A1(new_n844), .A2(new_n843), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n879), .A3(new_n846), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n837), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n883), .B1(new_n905), .B2(new_n880), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n888), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n443), .B(KEYINPUT57), .Z(new_n908));
  OAI21_X1  g722(.A(new_n701), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n894), .A2(new_n776), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(G54));
  NAND2_X1  g725(.A1(new_n905), .A2(new_n880), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n563), .A2(new_n557), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT120), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n901), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G60));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n630), .A2(new_n631), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n836), .A2(new_n840), .A3(new_n837), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n840), .B1(new_n836), .B2(new_n837), .ZN(new_n922));
  AND4_X1   g736(.A1(KEYINPUT53), .A2(new_n903), .A3(new_n879), .A4(new_n846), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n884), .B1(new_n924), .B2(new_n883), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n628), .B(KEYINPUT59), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n920), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n630), .B2(new_n631), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n888), .B2(new_n906), .ZN(new_n930));
  INV_X1    g744(.A(new_n901), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n919), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n889), .A2(new_n926), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n934), .B(KEYINPUT121), .C1(new_n935), .C2(new_n920), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(G63));
  XOR2_X1   g751(.A(new_n378), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n912), .A2(new_n653), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n912), .A2(new_n938), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n931), .B(new_n939), .C1(new_n940), .C2(new_n385), .ZN(new_n941));
  NAND2_X1  g755(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n942));
  OR2_X1    g756(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n941), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(G66));
  INV_X1    g760(.A(G224), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n515), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n824), .B2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n503), .B1(G898), .B2(new_n369), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G69));
  NOR2_X1   g765(.A1(new_n626), .A2(new_n673), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n782), .A2(new_n748), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n764), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(new_n787), .A3(new_n754), .A4(new_n783), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n695), .A2(new_n826), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n369), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(G900), .B2(new_n369), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT125), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n959), .B(new_n962), .C1(G900), .C2(new_n369), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n288), .B1(new_n295), .B2(new_n297), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n555), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n958), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n687), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n787), .A2(new_n783), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n756), .A2(new_n757), .A3(new_n623), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n743), .B(new_n676), .C1(new_n634), .C2(new_n664), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n970), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n966), .A2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n426), .B2(new_n665), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n976), .A2(new_n977), .B1(KEYINPUT126), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(KEYINPUT126), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  INV_X1    g798(.A(new_n824), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n298), .A2(new_n261), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT127), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n260), .A3(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n956), .A2(new_n985), .A3(new_n958), .ZN(new_n990));
  INV_X1    g804(.A(new_n984), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n988), .A2(new_n260), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n901), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n299), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n991), .B1(new_n996), .B2(new_n325), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n995), .B1(new_n848), .B2(new_n997), .ZN(G57));
endmodule


