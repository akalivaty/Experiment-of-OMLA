

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735;

  NOR2_X1 U373 ( .A1(G953), .A2(G237), .ZN(n496) );
  INV_X1 U374 ( .A(G953), .ZN(n724) );
  BUF_X1 U375 ( .A(n418), .Z(n702) );
  XNOR2_X1 U376 ( .A(n572), .B(KEYINPUT83), .ZN(n578) );
  NAND2_X1 U377 ( .A1(n678), .A2(n580), .ZN(n581) );
  INV_X2 U378 ( .A(G137), .ZN(n380) );
  NOR2_X1 U379 ( .A1(n647), .A2(G953), .ZN(n649) );
  NAND2_X1 U380 ( .A1(n351), .A2(n352), .ZN(n409) );
  NOR2_X1 U381 ( .A1(n403), .A2(n544), .ZN(n402) );
  XNOR2_X1 U382 ( .A(n575), .B(KEYINPUT40), .ZN(n733) );
  NOR2_X1 U383 ( .A1(n604), .A2(n585), .ZN(n684) );
  XNOR2_X1 U384 ( .A(n411), .B(KEYINPUT113), .ZN(n631) );
  XNOR2_X1 U385 ( .A(n373), .B(n353), .ZN(n565) );
  INV_X1 U386 ( .A(KEYINPUT94), .ZN(n363) );
  OR2_X1 U387 ( .A1(n695), .A2(G902), .ZN(n373) );
  NOR2_X1 U388 ( .A1(n601), .A2(n600), .ZN(n394) );
  INV_X1 U389 ( .A(n631), .ZN(n595) );
  AND2_X1 U390 ( .A1(n545), .A2(n415), .ZN(n544) );
  XNOR2_X1 U391 ( .A(n424), .B(n423), .ZN(n510) );
  XNOR2_X1 U392 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n423) );
  XNOR2_X1 U393 ( .A(G146), .B(G125), .ZN(n463) );
  XNOR2_X1 U394 ( .A(KEYINPUT3), .B(G119), .ZN(n456) );
  XNOR2_X1 U395 ( .A(n389), .B(n361), .ZN(n610) );
  XNOR2_X1 U396 ( .A(n611), .B(KEYINPUT92), .ZN(n723) );
  XNOR2_X1 U397 ( .A(n426), .B(n397), .ZN(n396) );
  XNOR2_X1 U398 ( .A(n422), .B(n398), .ZN(n397) );
  XNOR2_X1 U399 ( .A(n439), .B(n425), .ZN(n426) );
  XNOR2_X1 U400 ( .A(G128), .B(KEYINPUT103), .ZN(n422) );
  NAND2_X1 U401 ( .A1(n510), .A2(G221), .ZN(n395) );
  XNOR2_X1 U402 ( .A(n410), .B(KEYINPUT109), .ZN(n507) );
  INV_X1 U403 ( .A(KEYINPUT111), .ZN(n410) );
  XNOR2_X1 U404 ( .A(KEYINPUT110), .B(KEYINPUT9), .ZN(n506) );
  XNOR2_X1 U405 ( .A(G116), .B(G122), .ZN(n504) );
  XNOR2_X1 U406 ( .A(n437), .B(G128), .ZN(n512) );
  XNOR2_X1 U407 ( .A(G134), .B(G143), .ZN(n437) );
  XNOR2_X1 U408 ( .A(G113), .B(G143), .ZN(n490) );
  XOR2_X1 U409 ( .A(G104), .B(G122), .Z(n491) );
  XNOR2_X1 U410 ( .A(G131), .B(KEYINPUT12), .ZN(n492) );
  XOR2_X1 U411 ( .A(G140), .B(KEYINPUT11), .Z(n493) );
  XNOR2_X1 U412 ( .A(n463), .B(KEYINPUT10), .ZN(n722) );
  AND2_X1 U413 ( .A1(n369), .A2(n513), .ZN(n368) );
  XNOR2_X1 U414 ( .A(n565), .B(n359), .ZN(n616) );
  XNOR2_X1 U415 ( .A(n579), .B(KEYINPUT115), .ZN(n386) );
  XNOR2_X1 U416 ( .A(n391), .B(n362), .ZN(n390) );
  OR2_X1 U417 ( .A1(n678), .A2(n681), .ZN(n411) );
  XNOR2_X1 U418 ( .A(KEYINPUT15), .B(G902), .ZN(n652) );
  XOR2_X1 U419 ( .A(KEYINPUT82), .B(KEYINPUT105), .Z(n447) );
  XNOR2_X1 U420 ( .A(G137), .B(G146), .ZN(n448) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT106), .Z(n449) );
  XNOR2_X1 U422 ( .A(G119), .B(G110), .ZN(n425) );
  XNOR2_X1 U423 ( .A(KEYINPUT102), .B(KEYINPUT24), .ZN(n398) );
  XNOR2_X1 U424 ( .A(n512), .B(n438), .ZN(n453) );
  XNOR2_X1 U425 ( .A(KEYINPUT4), .B(G131), .ZN(n438) );
  NAND2_X1 U426 ( .A1(G234), .A2(G237), .ZN(n480) );
  INV_X1 U427 ( .A(G237), .ZN(n474) );
  INV_X1 U428 ( .A(G902), .ZN(n475) );
  XNOR2_X1 U429 ( .A(n374), .B(G107), .ZN(n713) );
  XNOR2_X1 U430 ( .A(G104), .B(G110), .ZN(n374) );
  XOR2_X1 U431 ( .A(G101), .B(G146), .Z(n442) );
  XOR2_X1 U432 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n465) );
  XNOR2_X1 U433 ( .A(n417), .B(n463), .ZN(n467) );
  XNOR2_X1 U434 ( .A(n399), .B(G143), .ZN(n417) );
  XNOR2_X1 U435 ( .A(KEYINPUT16), .B(G122), .ZN(n471) );
  NOR2_X1 U436 ( .A1(n723), .A2(KEYINPUT2), .ZN(n378) );
  NOR2_X1 U437 ( .A1(n629), .A2(n630), .ZN(n553) );
  AND2_X1 U438 ( .A1(n529), .A2(n622), .ZN(n624) );
  NOR2_X1 U439 ( .A1(n570), .A2(n569), .ZN(n365) );
  INV_X1 U440 ( .A(n616), .ZN(n604) );
  XNOR2_X1 U441 ( .A(n429), .B(n428), .ZN(n704) );
  XNOR2_X1 U442 ( .A(n722), .B(n427), .ZN(n428) );
  XNOR2_X1 U443 ( .A(n396), .B(n395), .ZN(n429) );
  XNOR2_X1 U444 ( .A(n413), .B(n412), .ZN(n699) );
  XNOR2_X1 U445 ( .A(n508), .B(n512), .ZN(n412) );
  XNOR2_X1 U446 ( .A(n511), .B(n509), .ZN(n413) );
  XNOR2_X1 U447 ( .A(n499), .B(n498), .ZN(n662) );
  XNOR2_X1 U448 ( .A(n722), .B(n497), .ZN(n498) );
  AND2_X1 U449 ( .A1(n658), .A2(G953), .ZN(n706) );
  XNOR2_X1 U450 ( .A(n384), .B(KEYINPUT91), .ZN(n646) );
  NAND2_X1 U451 ( .A1(n408), .A2(n376), .ZN(n384) );
  NAND2_X1 U452 ( .A1(n351), .A2(KEYINPUT2), .ZN(n408) );
  INV_X1 U453 ( .A(n388), .ZN(n376) );
  NAND2_X1 U454 ( .A1(n367), .A2(n366), .ZN(n514) );
  AND2_X1 U455 ( .A1(n370), .A2(n368), .ZN(n367) );
  XNOR2_X1 U456 ( .A(n524), .B(KEYINPUT32), .ZN(n406) );
  NOR2_X1 U457 ( .A1(n356), .A2(n580), .ZN(n414) );
  INV_X1 U458 ( .A(G143), .ZN(n385) );
  OR2_X1 U459 ( .A1(n707), .A2(n611), .ZN(n351) );
  AND2_X1 U460 ( .A1(n653), .A2(KEYINPUT2), .ZN(n352) );
  XOR2_X1 U461 ( .A(KEYINPUT73), .B(G469), .Z(n353) );
  OR2_X1 U462 ( .A1(n699), .A2(G902), .ZN(n354) );
  AND2_X1 U463 ( .A1(n476), .A2(G210), .ZN(n355) );
  XNOR2_X1 U464 ( .A(n462), .B(n461), .ZN(n634) );
  NAND2_X1 U465 ( .A1(n616), .A2(n612), .ZN(n356) );
  XNOR2_X1 U466 ( .A(n400), .B(n551), .ZN(n707) );
  INV_X1 U467 ( .A(n707), .ZN(n379) );
  NAND2_X1 U468 ( .A1(n485), .A2(n554), .ZN(n357) );
  XOR2_X1 U469 ( .A(n520), .B(KEYINPUT22), .Z(n358) );
  XOR2_X1 U470 ( .A(KEYINPUT67), .B(KEYINPUT1), .Z(n359) );
  XOR2_X1 U471 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n360) );
  XOR2_X1 U472 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n361) );
  XOR2_X1 U473 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n362) );
  XNOR2_X2 U474 ( .A(n536), .B(KEYINPUT112), .ZN(n678) );
  NOR2_X1 U475 ( .A1(n662), .A2(G902), .ZN(n501) );
  AND2_X2 U476 ( .A1(n378), .A2(n379), .ZN(n388) );
  XNOR2_X2 U477 ( .A(n364), .B(n363), .ZN(n545) );
  NAND2_X1 U478 ( .A1(n406), .A2(n405), .ZN(n364) );
  NAND2_X1 U479 ( .A1(n571), .A2(n365), .ZN(n572) );
  NAND2_X1 U480 ( .A1(n634), .A2(n489), .ZN(n366) );
  NAND2_X1 U481 ( .A1(n487), .A2(n489), .ZN(n369) );
  NAND2_X1 U482 ( .A1(n372), .A2(n371), .ZN(n370) );
  NOR2_X1 U483 ( .A1(n487), .A2(n489), .ZN(n371) );
  INV_X1 U484 ( .A(n634), .ZN(n372) );
  XNOR2_X1 U485 ( .A(n583), .B(n360), .ZN(n407) );
  XNOR2_X2 U486 ( .A(n375), .B(KEYINPUT95), .ZN(n583) );
  NAND2_X2 U487 ( .A1(n479), .A2(n478), .ZN(n375) );
  XNOR2_X2 U488 ( .A(n416), .B(n355), .ZN(n479) );
  NAND2_X1 U489 ( .A1(n377), .A2(n522), .ZN(n538) );
  NAND2_X1 U490 ( .A1(n377), .A2(n414), .ZN(n524) );
  AND2_X1 U491 ( .A1(n377), .A2(n527), .ZN(n650) );
  XNOR2_X2 U492 ( .A(n521), .B(n358), .ZN(n377) );
  XNOR2_X2 U493 ( .A(n380), .B(G140), .ZN(n439) );
  XNOR2_X2 U494 ( .A(n381), .B(KEYINPUT87), .ZN(n676) );
  NAND2_X1 U495 ( .A1(n382), .A2(n407), .ZN(n381) );
  INV_X1 U496 ( .A(n586), .ZN(n382) );
  NAND2_X1 U497 ( .A1(n564), .A2(n565), .ZN(n586) );
  NAND2_X1 U498 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X2 U499 ( .A(n383), .B(n486), .ZN(n519) );
  NAND2_X1 U500 ( .A1(n407), .A2(n357), .ZN(n383) );
  XNOR2_X1 U501 ( .A(n386), .B(n385), .ZN(G45) );
  XNOR2_X1 U502 ( .A(n386), .B(KEYINPUT89), .ZN(n591) );
  NAND2_X2 U503 ( .A1(n387), .A2(n409), .ZN(n418) );
  NAND2_X1 U504 ( .A1(n388), .A2(n653), .ZN(n387) );
  NAND2_X1 U505 ( .A1(n392), .A2(n390), .ZN(n389) );
  NAND2_X1 U506 ( .A1(n733), .A2(n735), .ZN(n391) );
  XNOR2_X1 U507 ( .A(n394), .B(n393), .ZN(n392) );
  INV_X1 U508 ( .A(KEYINPUT71), .ZN(n393) );
  XNOR2_X2 U509 ( .A(G128), .B(KEYINPUT4), .ZN(n399) );
  NAND2_X1 U510 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U511 ( .A1(n404), .A2(n550), .ZN(n401) );
  NAND2_X1 U512 ( .A1(n543), .A2(n542), .ZN(n403) );
  NAND2_X1 U513 ( .A1(n547), .A2(n548), .ZN(n404) );
  INV_X1 U514 ( .A(n650), .ZN(n405) );
  XNOR2_X1 U515 ( .A(n406), .B(G119), .ZN(G21) );
  XNOR2_X1 U516 ( .A(n721), .B(n444), .ZN(n695) );
  NOR2_X1 U517 ( .A1(n732), .A2(KEYINPUT44), .ZN(n415) );
  INV_X1 U518 ( .A(n479), .ZN(n552) );
  NAND2_X1 U519 ( .A1(n687), .A2(n652), .ZN(n416) );
  XNOR2_X1 U520 ( .A(n473), .B(n715), .ZN(n687) );
  XNOR2_X1 U521 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U522 ( .A(n597), .B(KEYINPUT80), .ZN(n598) );
  XNOR2_X1 U523 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U524 ( .A(KEYINPUT97), .B(KEYINPUT33), .ZN(n461) );
  XNOR2_X1 U525 ( .A(n453), .B(n452), .ZN(n458) );
  XNOR2_X1 U526 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n427) );
  XNOR2_X1 U527 ( .A(n468), .B(n443), .ZN(n444) );
  XNOR2_X1 U528 ( .A(n488), .B(KEYINPUT78), .ZN(n489) );
  NAND2_X1 U529 ( .A1(G234), .A2(n652), .ZN(n419) );
  XNOR2_X1 U530 ( .A(KEYINPUT20), .B(n419), .ZN(n430) );
  NAND2_X1 U531 ( .A1(n430), .A2(G221), .ZN(n420) );
  XNOR2_X1 U532 ( .A(n420), .B(KEYINPUT21), .ZN(n613) );
  INV_X1 U533 ( .A(KEYINPUT104), .ZN(n421) );
  XNOR2_X1 U534 ( .A(n613), .B(n421), .ZN(n516) );
  NAND2_X1 U535 ( .A1(n724), .A2(G234), .ZN(n424) );
  NOR2_X1 U536 ( .A1(n704), .A2(G902), .ZN(n434) );
  NAND2_X1 U537 ( .A1(n430), .A2(G217), .ZN(n432) );
  XNOR2_X1 U538 ( .A(KEYINPUT85), .B(KEYINPUT25), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U540 ( .A(n434), .B(n433), .ZN(n560) );
  INV_X1 U541 ( .A(n560), .ZN(n523) );
  NAND2_X1 U542 ( .A1(n516), .A2(n523), .ZN(n436) );
  INV_X1 U543 ( .A(KEYINPUT68), .ZN(n435) );
  XNOR2_X2 U544 ( .A(n436), .B(n435), .ZN(n617) );
  XNOR2_X1 U545 ( .A(n439), .B(n453), .ZN(n721) );
  XNOR2_X1 U546 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n713), .B(n440), .ZN(n468) );
  NAND2_X1 U548 ( .A1(G227), .A2(n724), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U550 ( .A1(n617), .A2(n616), .ZN(n445) );
  XNOR2_X1 U551 ( .A(n445), .B(KEYINPUT81), .ZN(n529) );
  NAND2_X1 U552 ( .A1(n496), .A2(G210), .ZN(n446) );
  XNOR2_X1 U553 ( .A(n447), .B(n446), .ZN(n451) );
  XNOR2_X1 U554 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U555 ( .A(G116), .B(G113), .ZN(n455) );
  XNOR2_X1 U556 ( .A(G101), .B(KEYINPUT74), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n457) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n470) );
  XNOR2_X1 U559 ( .A(n458), .B(n470), .ZN(n655) );
  NAND2_X1 U560 ( .A1(n655), .A2(n475), .ZN(n460) );
  INV_X1 U561 ( .A(G472), .ZN(n459) );
  XNOR2_X1 U562 ( .A(n460), .B(n459), .ZN(n567) );
  XNOR2_X1 U563 ( .A(n567), .B(KEYINPUT6), .ZN(n580) );
  NAND2_X1 U564 ( .A1(n529), .A2(n580), .ZN(n462) );
  NAND2_X1 U565 ( .A1(G224), .A2(n724), .ZN(n464) );
  XNOR2_X1 U566 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n469), .B(n468), .ZN(n473) );
  INV_X1 U569 ( .A(n470), .ZN(n472) );
  XNOR2_X1 U570 ( .A(n472), .B(n471), .ZN(n715) );
  NAND2_X1 U571 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U572 ( .A1(n476), .A2(G214), .ZN(n477) );
  XNOR2_X1 U573 ( .A(n477), .B(KEYINPUT99), .ZN(n606) );
  INV_X1 U574 ( .A(n606), .ZN(n478) );
  XNOR2_X1 U575 ( .A(n480), .B(KEYINPUT14), .ZN(n482) );
  NAND2_X1 U576 ( .A1(n482), .A2(G902), .ZN(n481) );
  XNOR2_X1 U577 ( .A(n481), .B(KEYINPUT101), .ZN(n555) );
  NOR2_X1 U578 ( .A1(G898), .A2(n724), .ZN(n717) );
  NAND2_X1 U579 ( .A1(n555), .A2(n717), .ZN(n485) );
  NAND2_X1 U580 ( .A1(G952), .A2(n482), .ZN(n641) );
  NOR2_X1 U581 ( .A1(n641), .A2(G953), .ZN(n484) );
  INV_X1 U582 ( .A(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U583 ( .A(n484), .B(n483), .ZN(n554) );
  INV_X1 U584 ( .A(KEYINPUT0), .ZN(n486) );
  INV_X1 U585 ( .A(n519), .ZN(n487) );
  XNOR2_X1 U586 ( .A(KEYINPUT34), .B(KEYINPUT86), .ZN(n488) );
  XNOR2_X1 U587 ( .A(n491), .B(n490), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U589 ( .A(n495), .B(n494), .Z(n499) );
  NAND2_X1 U590 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT13), .ZN(n500) );
  XNOR2_X1 U592 ( .A(n501), .B(n500), .ZN(n503) );
  INV_X1 U593 ( .A(G475), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n503), .B(n502), .ZN(n535) );
  XOR2_X1 U595 ( .A(KEYINPUT7), .B(G107), .Z(n505) );
  XNOR2_X1 U596 ( .A(n505), .B(n504), .ZN(n509) );
  XNOR2_X1 U597 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U598 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U599 ( .A(G478), .B(n354), .ZN(n534) );
  INV_X1 U600 ( .A(n534), .ZN(n515) );
  OR2_X1 U601 ( .A1(n535), .A2(n515), .ZN(n576) );
  INV_X1 U602 ( .A(n576), .ZN(n513) );
  XNOR2_X2 U603 ( .A(n514), .B(KEYINPUT35), .ZN(n732) );
  INV_X1 U604 ( .A(KEYINPUT44), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n535), .A2(n515), .ZN(n629) );
  INV_X1 U606 ( .A(n516), .ZN(n517) );
  NOR2_X1 U607 ( .A1(n629), .A2(n517), .ZN(n518) );
  INV_X1 U608 ( .A(KEYINPUT79), .ZN(n520) );
  INV_X1 U609 ( .A(n580), .ZN(n522) );
  INV_X1 U610 ( .A(n523), .ZN(n525) );
  XNOR2_X1 U611 ( .A(n525), .B(KEYINPUT114), .ZN(n612) );
  AND2_X1 U612 ( .A1(n525), .A2(n567), .ZN(n526) );
  AND2_X1 U613 ( .A1(n604), .A2(n526), .ZN(n527) );
  INV_X1 U614 ( .A(KEYINPUT66), .ZN(n528) );
  NAND2_X1 U615 ( .A1(n545), .A2(n528), .ZN(n543) );
  INV_X1 U616 ( .A(n567), .ZN(n622) );
  NAND2_X1 U617 ( .A1(n624), .A2(n519), .ZN(n530) );
  XNOR2_X1 U618 ( .A(n530), .B(KEYINPUT31), .ZN(n682) );
  NAND2_X1 U619 ( .A1(n565), .A2(n617), .ZN(n570) );
  NOR2_X1 U620 ( .A1(n570), .A2(n622), .ZN(n531) );
  AND2_X1 U621 ( .A1(n519), .A2(n531), .ZN(n669) );
  OR2_X1 U622 ( .A1(n682), .A2(n669), .ZN(n533) );
  INV_X1 U623 ( .A(KEYINPUT107), .ZN(n532) );
  XNOR2_X1 U624 ( .A(n533), .B(n532), .ZN(n537) );
  AND2_X1 U625 ( .A1(n534), .A2(n535), .ZN(n681) );
  NOR2_X1 U626 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U627 ( .A1(n537), .A2(n595), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n538), .B(KEYINPUT93), .ZN(n540) );
  NOR2_X1 U629 ( .A1(n616), .A2(n612), .ZN(n539) );
  NAND2_X1 U630 ( .A1(n540), .A2(n539), .ZN(n667) );
  AND2_X1 U631 ( .A1(n541), .A2(n667), .ZN(n542) );
  NOR2_X1 U632 ( .A1(n732), .A2(n549), .ZN(n548) );
  INV_X1 U633 ( .A(n545), .ZN(n546) );
  NAND2_X1 U634 ( .A1(n546), .A2(KEYINPUT66), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n549), .A2(KEYINPUT66), .ZN(n550) );
  XNOR2_X1 U636 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n551) );
  XNOR2_X1 U637 ( .A(n552), .B(KEYINPUT38), .ZN(n627) );
  NAND2_X1 U638 ( .A1(n627), .A2(n478), .ZN(n630) );
  XNOR2_X1 U639 ( .A(n553), .B(KEYINPUT41), .ZN(n642) );
  XNOR2_X1 U640 ( .A(KEYINPUT28), .B(KEYINPUT116), .ZN(n563) );
  INV_X1 U641 ( .A(n554), .ZN(n558) );
  NAND2_X1 U642 ( .A1(n555), .A2(G953), .ZN(n556) );
  NOR2_X1 U643 ( .A1(G900), .A2(n556), .ZN(n557) );
  NOR2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n569) );
  NOR2_X1 U645 ( .A1(n613), .A2(n569), .ZN(n559) );
  XNOR2_X1 U646 ( .A(KEYINPUT72), .B(n559), .ZN(n561) );
  NAND2_X1 U647 ( .A1(n561), .A2(n525), .ZN(n582) );
  NOR2_X1 U648 ( .A1(n582), .A2(n567), .ZN(n562) );
  XNOR2_X1 U649 ( .A(n563), .B(n562), .ZN(n564) );
  NOR2_X1 U650 ( .A1(n642), .A2(n586), .ZN(n566) );
  XOR2_X1 U651 ( .A(KEYINPUT42), .B(n566), .Z(n735) );
  NOR2_X1 U652 ( .A1(n606), .A2(n567), .ZN(n568) );
  XNOR2_X1 U653 ( .A(KEYINPUT30), .B(n568), .ZN(n571) );
  NAND2_X1 U654 ( .A1(n578), .A2(n627), .ZN(n574) );
  XOR2_X1 U655 ( .A(KEYINPUT77), .B(KEYINPUT39), .Z(n573) );
  XNOR2_X1 U656 ( .A(n574), .B(n573), .ZN(n602) );
  NAND2_X1 U657 ( .A1(n602), .A2(n678), .ZN(n575) );
  NOR2_X1 U658 ( .A1(n576), .A2(n552), .ZN(n577) );
  NAND2_X1 U659 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n603) );
  NAND2_X1 U661 ( .A1(n603), .A2(n583), .ZN(n584) );
  XNOR2_X1 U662 ( .A(n584), .B(KEYINPUT36), .ZN(n585) );
  INV_X1 U663 ( .A(KEYINPUT47), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n587), .A2(n676), .ZN(n588) );
  NOR2_X1 U665 ( .A1(KEYINPUT88), .A2(n588), .ZN(n589) );
  NOR2_X1 U666 ( .A1(n684), .A2(n589), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n601) );
  INV_X1 U668 ( .A(n676), .ZN(n592) );
  NAND2_X1 U669 ( .A1(KEYINPUT88), .A2(n592), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n593), .A2(n595), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n594), .A2(KEYINPUT47), .ZN(n599) );
  NOR2_X1 U672 ( .A1(n631), .A2(KEYINPUT47), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n676), .A2(n596), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n602), .A2(n681), .ZN(n686) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U678 ( .A(n607), .B(KEYINPUT43), .Z(n608) );
  NAND2_X1 U679 ( .A1(n608), .A2(n552), .ZN(n651) );
  AND2_X1 U680 ( .A1(n686), .A2(n651), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n615) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(n620) );
  NOR2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U686 ( .A(KEYINPUT50), .B(n618), .Z(n619) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U688 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U689 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U690 ( .A(KEYINPUT51), .B(n625), .Z(n626) );
  NOR2_X1 U691 ( .A1(n642), .A2(n626), .ZN(n637) );
  NOR2_X1 U692 ( .A1(n627), .A2(n478), .ZN(n628) );
  NOR2_X1 U693 ( .A1(n629), .A2(n628), .ZN(n633) );
  NOR2_X1 U694 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U695 ( .A1(n633), .A2(n632), .ZN(n635) );
  NOR2_X1 U696 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U697 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U698 ( .A(n638), .B(KEYINPUT121), .Z(n639) );
  XNOR2_X1 U699 ( .A(KEYINPUT52), .B(n639), .ZN(n640) );
  NOR2_X1 U700 ( .A1(n641), .A2(n640), .ZN(n644) );
  NOR2_X1 U701 ( .A1(n634), .A2(n642), .ZN(n643) );
  NOR2_X1 U702 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U703 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U704 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n648) );
  XNOR2_X1 U705 ( .A(n649), .B(n648), .ZN(G75) );
  XOR2_X1 U706 ( .A(G110), .B(n650), .Z(G12) );
  XNOR2_X1 U707 ( .A(n651), .B(G140), .ZN(G42) );
  INV_X1 U708 ( .A(n652), .ZN(n653) );
  NAND2_X1 U709 ( .A1(n418), .A2(G472), .ZN(n657) );
  XOR2_X1 U710 ( .A(KEYINPUT98), .B(KEYINPUT62), .Z(n654) );
  XNOR2_X1 U711 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U712 ( .A(n657), .B(n656), .ZN(n659) );
  INV_X1 U713 ( .A(G952), .ZN(n658) );
  NOR2_X2 U714 ( .A1(n659), .A2(n706), .ZN(n661) );
  XNOR2_X1 U715 ( .A(KEYINPUT117), .B(KEYINPUT63), .ZN(n660) );
  XNOR2_X1 U716 ( .A(n661), .B(n660), .ZN(G57) );
  NAND2_X1 U717 ( .A1(n418), .A2(G475), .ZN(n664) );
  XOR2_X1 U718 ( .A(n662), .B(KEYINPUT59), .Z(n663) );
  XNOR2_X1 U719 ( .A(n664), .B(n663), .ZN(n665) );
  NOR2_X2 U720 ( .A1(n665), .A2(n706), .ZN(n666) );
  XNOR2_X1 U721 ( .A(n666), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U722 ( .A(G101), .B(n667), .ZN(G3) );
  NAND2_X1 U723 ( .A1(n678), .A2(n669), .ZN(n668) );
  XNOR2_X1 U724 ( .A(n668), .B(G104), .ZN(G6) );
  XNOR2_X1 U725 ( .A(G107), .B(KEYINPUT118), .ZN(n673) );
  XOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n671) );
  NAND2_X1 U727 ( .A1(n669), .A2(n681), .ZN(n670) );
  XNOR2_X1 U728 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U729 ( .A(n673), .B(n672), .ZN(G9) );
  XOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U731 ( .A1(n676), .A2(n681), .ZN(n674) );
  XNOR2_X1 U732 ( .A(n675), .B(n674), .ZN(G30) );
  NAND2_X1 U733 ( .A1(n678), .A2(n676), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n677), .B(G146), .ZN(G48) );
  XOR2_X1 U735 ( .A(G113), .B(KEYINPUT119), .Z(n680) );
  NAND2_X1 U736 ( .A1(n682), .A2(n678), .ZN(n679) );
  XNOR2_X1 U737 ( .A(n680), .B(n679), .ZN(G15) );
  NAND2_X1 U738 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U739 ( .A(n683), .B(G116), .ZN(G18) );
  XNOR2_X1 U740 ( .A(G125), .B(n684), .ZN(n685) );
  XNOR2_X1 U741 ( .A(n685), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U742 ( .A(G134), .B(n686), .ZN(G36) );
  NAND2_X1 U743 ( .A1(n418), .A2(G210), .ZN(n691) );
  XNOR2_X1 U744 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n688) );
  XNOR2_X1 U745 ( .A(n688), .B(KEYINPUT96), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n687), .B(n689), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X2 U748 ( .A1(n692), .A2(n706), .ZN(n693) );
  XNOR2_X1 U749 ( .A(n693), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U750 ( .A1(n702), .A2(G469), .ZN(n697) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U752 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n706), .A2(n698), .ZN(G54) );
  NAND2_X1 U754 ( .A1(n702), .A2(G478), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U756 ( .A1(n706), .A2(n701), .ZN(G63) );
  NAND2_X1 U757 ( .A1(n702), .A2(G217), .ZN(n703) );
  XNOR2_X1 U758 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U760 ( .A1(n379), .A2(n724), .ZN(n712) );
  XOR2_X1 U761 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n709) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U764 ( .A1(n710), .A2(G898), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n719) );
  XOR2_X1 U766 ( .A(n713), .B(KEYINPUT124), .Z(n714) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U769 ( .A(n719), .B(n718), .Z(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT125), .B(n720), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n726) );
  XNOR2_X1 U772 ( .A(n723), .B(n726), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U774 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U776 ( .A1(G953), .A2(n728), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U778 ( .A(KEYINPUT126), .B(n731), .ZN(G72) );
  XOR2_X1 U779 ( .A(G122), .B(n732), .Z(G24) );
  XOR2_X1 U780 ( .A(G131), .B(n733), .Z(n734) );
  XNOR2_X1 U781 ( .A(KEYINPUT127), .B(n734), .ZN(G33) );
  XNOR2_X1 U782 ( .A(n735), .B(G137), .ZN(G39) );
endmodule

