

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  NOR2_X1 U319 ( .A1(n471), .A2(n470), .ZN(n485) );
  XNOR2_X1 U320 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U321 ( .A(n488), .B(KEYINPUT96), .ZN(n489) );
  XNOR2_X1 U322 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U323 ( .A(n454), .B(KEYINPUT121), .ZN(n562) );
  XOR2_X1 U324 ( .A(n464), .B(KEYINPUT25), .Z(n287) );
  XOR2_X1 U325 ( .A(n399), .B(KEYINPUT84), .Z(n288) );
  XOR2_X1 U326 ( .A(n373), .B(KEYINPUT29), .Z(n289) );
  XOR2_X1 U327 ( .A(G29GAT), .B(G43GAT), .Z(n290) );
  NOR2_X1 U328 ( .A1(n387), .A2(n557), .ZN(n388) );
  AND2_X1 U329 ( .A1(n465), .A2(n287), .ZN(n466) );
  NOR2_X1 U330 ( .A1(n469), .A2(n531), .ZN(n462) );
  XNOR2_X1 U331 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n436) );
  XNOR2_X1 U332 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U333 ( .A(n437), .B(n436), .ZN(n453) );
  XNOR2_X1 U334 ( .A(n340), .B(n339), .ZN(n346) );
  XNOR2_X1 U335 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U336 ( .A(n490), .B(n489), .ZN(n515) );
  XOR2_X1 U337 ( .A(n363), .B(n362), .Z(n566) );
  XOR2_X1 U338 ( .A(n389), .B(KEYINPUT41), .Z(n552) );
  XOR2_X1 U339 ( .A(n452), .B(n451), .Z(n524) );
  XNOR2_X1 U340 ( .A(n492), .B(KEYINPUT38), .ZN(n501) );
  XNOR2_X1 U341 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n459) );
  XNOR2_X1 U342 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n292) );
  XNOR2_X1 U344 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n310) );
  XOR2_X1 U346 ( .A(G85GAT), .B(G127GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(G141GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U349 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n296) );
  XNOR2_X1 U350 ( .A(G148GAT), .B(G57GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(n298), .B(n297), .Z(n304) );
  XNOR2_X1 U353 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n299), .B(KEYINPUT2), .ZN(n423) );
  XOR2_X1 U355 ( .A(G162GAT), .B(n423), .Z(n301) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(n302), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n305), .B(KEYINPUT1), .Z(n308) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n306), .B(KEYINPUT0), .ZN(n449) );
  XNOR2_X1 U363 ( .A(G1GAT), .B(n449), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n517) );
  INV_X1 U366 ( .A(n517), .ZN(n467) );
  XOR2_X1 U367 ( .A(G78GAT), .B(G155GAT), .Z(n312) );
  XNOR2_X1 U368 ( .A(G22GAT), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n314) );
  XNOR2_X1 U371 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n447) );
  XOR2_X1 U374 ( .A(n447), .B(G71GAT), .Z(n316) );
  XOR2_X1 U375 ( .A(G1GAT), .B(G8GAT), .Z(n349) );
  XNOR2_X1 U376 ( .A(n349), .B(G183GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U378 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U379 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U381 ( .A(n321), .B(KEYINPUT81), .Z(n324) );
  XNOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n322), .B(KEYINPUT72), .ZN(n338) );
  XNOR2_X1 U384 ( .A(n338), .B(KEYINPUT12), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n486) );
  INV_X1 U387 ( .A(n486), .ZN(n574) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XOR2_X1 U389 ( .A(G99GAT), .B(G85GAT), .Z(n369) );
  XNOR2_X1 U390 ( .A(n450), .B(n369), .ZN(n328) );
  XOR2_X1 U391 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n333) );
  INV_X1 U393 ( .A(n333), .ZN(n332) );
  XOR2_X1 U394 ( .A(KEYINPUT73), .B(KEYINPUT76), .Z(n330) );
  XNOR2_X1 U395 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n329) );
  XNOR2_X1 U396 ( .A(n330), .B(n329), .ZN(n334) );
  INV_X1 U397 ( .A(n334), .ZN(n331) );
  NAND2_X1 U398 ( .A1(n332), .A2(n331), .ZN(n336) );
  NAND2_X1 U399 ( .A1(n334), .A2(n333), .ZN(n335) );
  NAND2_X1 U400 ( .A1(n336), .A2(n335), .ZN(n340) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n341), .B(G148GAT), .ZN(n422) );
  XOR2_X1 U404 ( .A(G92GAT), .B(KEYINPUT75), .Z(n343) );
  XNOR2_X1 U405 ( .A(G176GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U407 ( .A(G204GAT), .B(n344), .Z(n404) );
  XNOR2_X1 U408 ( .A(n422), .B(n404), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n389) );
  XOR2_X1 U410 ( .A(G15GAT), .B(G113GAT), .Z(n348) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G36GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U413 ( .A(n350), .B(n349), .Z(n355) );
  XNOR2_X1 U414 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n290), .B(n351), .ZN(n373) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n289), .B(n352), .ZN(n353) );
  XOR2_X1 U418 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XNOR2_X1 U419 ( .A(n353), .B(n431), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n357) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(G197GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U424 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n359) );
  XNOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT71), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  INV_X1 U428 ( .A(n566), .ZN(n559) );
  NAND2_X1 U429 ( .A1(n552), .A2(n559), .ZN(n366) );
  XOR2_X1 U430 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n364) );
  XNOR2_X1 U431 ( .A(KEYINPUT109), .B(n364), .ZN(n365) );
  XOR2_X1 U432 ( .A(n366), .B(n365), .Z(n367) );
  NOR2_X1 U433 ( .A1(n574), .A2(n367), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n368), .B(KEYINPUT111), .ZN(n387) );
  XOR2_X1 U435 ( .A(KEYINPUT79), .B(KEYINPUT9), .Z(n371) );
  XOR2_X1 U436 ( .A(G36GAT), .B(G190GAT), .Z(n401) );
  XNOR2_X1 U437 ( .A(n369), .B(n401), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U439 ( .A(n372), .B(KEYINPUT66), .Z(n378) );
  XOR2_X1 U440 ( .A(G50GAT), .B(G162GAT), .Z(n430) );
  XOR2_X1 U441 ( .A(n373), .B(n430), .Z(n375) );
  NAND2_X1 U442 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U444 ( .A(G218GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n380) );
  XNOR2_X1 U447 ( .A(KEYINPUT10), .B(KEYINPUT78), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U449 ( .A(KEYINPUT65), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(G134GAT), .B(G106GAT), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n472) );
  INV_X1 U454 ( .A(n472), .ZN(n557) );
  XNOR2_X1 U455 ( .A(n388), .B(KEYINPUT47), .ZN(n395) );
  XOR2_X1 U456 ( .A(KEYINPUT36), .B(n557), .Z(n578) );
  NOR2_X1 U457 ( .A1(n578), .A2(n486), .ZN(n390) );
  XOR2_X1 U458 ( .A(KEYINPUT45), .B(n390), .Z(n391) );
  NOR2_X1 U459 ( .A1(n389), .A2(n391), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n392), .B(KEYINPUT112), .ZN(n393) );
  NAND2_X1 U461 ( .A1(n393), .A2(n566), .ZN(n394) );
  NAND2_X1 U462 ( .A1(n395), .A2(n394), .ZN(n397) );
  INV_X1 U463 ( .A(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n547) );
  INV_X1 U465 ( .A(n547), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n398), .B(KEYINPUT19), .ZN(n399) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(G183GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n288), .B(n400), .ZN(n445) );
  XOR2_X1 U469 ( .A(n401), .B(KEYINPUT93), .Z(n403) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U472 ( .A(n405), .B(n404), .Z(n411) );
  XOR2_X1 U473 ( .A(KEYINPUT21), .B(G218GAT), .Z(n407) );
  XNOR2_X1 U474 ( .A(KEYINPUT87), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U476 ( .A(G197GAT), .B(n408), .Z(n434) );
  INV_X1 U477 ( .A(n434), .ZN(n409) );
  XOR2_X1 U478 ( .A(G8GAT), .B(n409), .Z(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n445), .B(n412), .ZN(n521) );
  XNOR2_X1 U481 ( .A(KEYINPUT117), .B(n521), .ZN(n413) );
  NAND2_X1 U482 ( .A1(n414), .A2(n413), .ZN(n417) );
  XNOR2_X1 U483 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n415) );
  XOR2_X1 U484 ( .A(n415), .B(KEYINPUT54), .Z(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n418) );
  NOR2_X1 U486 ( .A1(n467), .A2(n418), .ZN(n565) );
  XOR2_X1 U487 ( .A(KEYINPUT86), .B(KEYINPUT89), .Z(n420) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U490 ( .A(n421), .B(KEYINPUT88), .Z(n425) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U493 ( .A(G204GAT), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U494 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U496 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U499 ( .A(n435), .B(n434), .Z(n469) );
  NAND2_X1 U500 ( .A1(n565), .A2(n469), .ZN(n437) );
  XOR2_X1 U501 ( .A(KEYINPUT85), .B(G176GAT), .Z(n439) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U504 ( .A(n440), .B(KEYINPUT20), .Z(n444) );
  XOR2_X1 U505 ( .A(KEYINPUT83), .B(G99GAT), .Z(n442) );
  XNOR2_X1 U506 ( .A(G43GAT), .B(G190GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U508 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U510 ( .A(n524), .ZN(n531) );
  NAND2_X1 U511 ( .A1(n453), .A2(n531), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n562), .A2(n552), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n456) );
  XOR2_X1 U514 ( .A(G176GAT), .B(KEYINPUT123), .Z(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  NAND2_X1 U517 ( .A1(n557), .A2(n562), .ZN(n460) );
  NOR2_X1 U518 ( .A1(n389), .A2(n566), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT77), .B(n461), .Z(n491) );
  XOR2_X1 U520 ( .A(n462), .B(KEYINPUT26), .Z(n544) );
  XNOR2_X1 U521 ( .A(KEYINPUT27), .B(n521), .ZN(n468) );
  OR2_X1 U522 ( .A1(n544), .A2(n468), .ZN(n465) );
  OR2_X1 U523 ( .A1(n524), .A2(n521), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n469), .A2(n463), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n468), .A2(n517), .ZN(n545) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT28), .ZN(n527) );
  NAND2_X1 U528 ( .A1(n545), .A2(n527), .ZN(n533) );
  NOR2_X1 U529 ( .A1(n531), .A2(n533), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n574), .A2(n472), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(KEYINPUT82), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT16), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n485), .A2(n475), .ZN(n504) );
  NAND2_X1 U534 ( .A1(n491), .A2(n504), .ZN(n482) );
  NOR2_X1 U535 ( .A1(n517), .A2(n482), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(n476), .Z(n477) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U538 ( .A1(n521), .A2(n482), .ZN(n478) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n478), .Z(G1325GAT) );
  NOR2_X1 U540 ( .A1(n524), .A2(n482), .ZN(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT35), .B(KEYINPUT94), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n527), .A2(n482), .ZN(n484) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT95), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  NOR2_X1 U547 ( .A1(n485), .A2(n578), .ZN(n487) );
  NAND2_X1 U548 ( .A1(n487), .A2(n486), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT97), .B(KEYINPUT37), .Z(n488) );
  NAND2_X1 U550 ( .A1(n515), .A2(n491), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n501), .A2(n517), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT98), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n501), .A2(n521), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT99), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  NOR2_X1 U558 ( .A1(n501), .A2(n524), .ZN(n499) );
  XNOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U561 ( .A(G43GAT), .B(n500), .Z(G1330GAT) );
  NOR2_X1 U562 ( .A1(n501), .A2(n527), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  AND2_X1 U565 ( .A1(n566), .A2(n552), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n516), .A2(n504), .ZN(n511) );
  NOR2_X1 U567 ( .A1(n517), .A2(n511), .ZN(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n507), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n521), .A2(n511), .ZN(n508) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n524), .A2(n511), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT103), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n527), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n517), .A2(n526), .ZN(n519) );
  XNOR2_X1 U582 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n526), .ZN(n525) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n414), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n559), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U599 ( .A1(n541), .A2(n552), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n540) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n538) );
  NAND2_X1 U603 ( .A1(n541), .A2(n574), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U607 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  INV_X1 U609 ( .A(n544), .ZN(n564) );
  NAND2_X1 U610 ( .A1(n545), .A2(n564), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n559), .A2(n556), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(n551), .Z(n554) );
  NAND2_X1 U618 ( .A1(n556), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n556), .A2(n574), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n559), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n574), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n566), .A2(n577), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(KEYINPUT124), .B(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U637 ( .A(n577), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n575), .A2(n389), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

