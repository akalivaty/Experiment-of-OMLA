//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT72), .B(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT73), .B(G155gat), .Z(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(KEYINPUT2), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n215), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n216));
  XOR2_X1   g015(.A(G127gat), .B(G134gat), .Z(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n218), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G225gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n219), .B2(new_n222), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT5), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n233), .B(new_n220), .C1(new_n221), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n214), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n224), .A4(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n227), .A2(new_n231), .A3(new_n232), .A4(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n227), .A2(new_n231), .A3(new_n240), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT76), .B1(new_n240), .B2(KEYINPUT5), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G1gat), .B(G29gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT0), .ZN(new_n246));
  XNOR2_X1  g045(.A(G57gat), .B(G85gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(new_n247), .Z(new_n248));
  AOI21_X1  g047(.A(KEYINPUT6), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G64gat), .B(G92gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(G183gat), .B2(G190gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT65), .B(G169gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI221_X1 g071(.A(new_n266), .B1(new_n267), .B2(new_n269), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(new_n271), .B2(new_n261), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n267), .B(KEYINPUT66), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n266), .B(new_n276), .C1(new_n277), .C2(new_n269), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT27), .B(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT28), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT26), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n264), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n263), .A2(new_n284), .B1(new_n287), .B2(new_n281), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n283), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n260), .B1(new_n279), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT70), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OR3_X1    g093(.A1(new_n283), .A2(new_n286), .A3(new_n288), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n278), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G226gat), .A3(G233gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT69), .B(G211gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G218gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n304), .B2(KEYINPUT22), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n291), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n297), .A2(new_n292), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n259), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(new_n259), .A3(new_n312), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n256), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT31), .B(G50gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n321), .B(G22gat), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n221), .A2(new_n235), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n307), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n260), .A3(new_n221), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n233), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n325), .A2(new_n326), .ZN(new_n330));
  OAI211_X1 g129(.A(G228gat), .B(G233gat), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT77), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n221), .A2(new_n235), .B1(G228gat), .B2(G233gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n325), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n331), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n323), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n322), .A3(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n220), .B1(new_n279), .B2(new_n289), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n295), .A2(new_n218), .A3(new_n296), .ZN(new_n345));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n346), .B(KEYINPUT64), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT34), .Z(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n345), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n347), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G15gat), .B(G43gat), .Z(new_n355));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n348), .B1(new_n344), .B2(new_n345), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n354), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  AOI221_X4 g159(.A(new_n358), .B1(KEYINPUT33), .B2(new_n357), .C1(new_n351), .C2(new_n347), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n350), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n350), .A3(new_n362), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n349), .B(KEYINPUT34), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n357), .B1(new_n359), .B2(KEYINPUT33), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n359), .A2(new_n358), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n370), .B2(new_n361), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n343), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT35), .B1(new_n320), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n318), .A2(KEYINPUT35), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n251), .A2(KEYINPUT79), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n227), .A2(new_n240), .A3(new_n231), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(KEYINPUT76), .C1(KEYINPUT5), .C2(new_n240), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n250), .A4(new_n241), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n249), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n255), .ZN(new_n383));
  INV_X1    g182(.A(new_n366), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n363), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n376), .A2(new_n383), .A3(new_n385), .A4(new_n343), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n254), .B1(new_n251), .B2(new_n249), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n343), .A2(new_n388), .A3(new_n318), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n377), .A2(new_n381), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT39), .B1(new_n223), .B2(new_n225), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n225), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n225), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n394), .B(new_n248), .C1(KEYINPUT39), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT40), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n390), .A2(new_n318), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n313), .ZN(new_n401));
  INV_X1    g200(.A(new_n259), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT37), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT38), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT80), .B1(new_n299), .B2(new_n307), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n294), .A2(new_n298), .A3(new_n406), .A4(new_n310), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n309), .A2(new_n311), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n307), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT37), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n410), .B2(KEYINPUT37), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n404), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n316), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n308), .A2(new_n312), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT37), .ZN(new_n417));
  INV_X1    g216(.A(new_n403), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n313), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n419), .B2(KEYINPUT38), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n382), .A2(new_n414), .A3(new_n255), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n389), .B1(new_n422), .B2(new_n343), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT36), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n365), .B2(new_n372), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT36), .B1(new_n366), .B2(new_n371), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n387), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT83), .ZN(new_n431));
  XOR2_X1   g230(.A(G113gat), .B(G141gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G169gat), .B(G197gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n433), .A2(new_n435), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n431), .B(new_n432), .Z(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n434), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n436), .A3(KEYINPUT12), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT15), .ZN(new_n444));
  NOR2_X1   g243(.A1(G43gat), .A2(G50gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G43gat), .A2(G50gat), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G36gat), .ZN(new_n449));
  AND2_X1   g248(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G29gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  INV_X1    g255(.A(G50gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G43gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(KEYINPUT84), .A2(G50gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n448), .B1(new_n455), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n447), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT15), .B1(new_n465), .B2(new_n445), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n452), .B2(new_n454), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(G1gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT16), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(G1gat), .ZN(new_n473));
  OAI21_X1  g272(.A(G8gat), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G15gat), .B(G22gat), .Z(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n470), .ZN(new_n476));
  INV_X1    g275(.A(G8gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n471), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n468), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n482), .B(KEYINPUT13), .Z(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n482), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT17), .B1(new_n464), .B2(new_n467), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n472), .A2(new_n473), .A3(G8gat), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT17), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n455), .A2(new_n448), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n452), .A2(new_n454), .B1(new_n461), .B2(new_n462), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n490), .B(new_n491), .C1(new_n492), .C2(new_n448), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n486), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT85), .B1(new_n468), .B2(new_n480), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT85), .A4(new_n493), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n485), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n484), .B1(new_n498), .B2(KEYINPUT18), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT18), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n500), .B(new_n485), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n443), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n499), .A2(new_n501), .ZN(new_n504));
  INV_X1    g303(.A(new_n443), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR4_X1   g305(.A1(new_n499), .A2(new_n443), .A3(new_n501), .A4(KEYINPUT86), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n428), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515));
  INV_X1    g314(.A(G85gat), .ZN(new_n516));
  INV_X1    g315(.A(G92gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(KEYINPUT8), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n522));
  AND2_X1   g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(KEYINPUT91), .B(new_n521), .C1(new_n516), .C2(new_n517), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n524), .A2(KEYINPUT92), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT92), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G99gat), .B(G106gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n529), .B(new_n518), .C1(new_n526), .C2(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT93), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n526), .A2(new_n527), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n529), .A4(new_n518), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n468), .ZN(new_n538));
  AND2_X1   g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n486), .A2(new_n493), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n533), .A3(new_n536), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n542), .A2(new_n533), .A3(KEYINPUT94), .A4(new_n536), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT95), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n546), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n537), .A2(new_n468), .B1(KEYINPUT41), .B2(new_n539), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n548), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(KEYINPUT96), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT96), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n554), .B1(new_n553), .B2(new_n548), .ZN(new_n558));
  AOI211_X1 g357(.A(KEYINPUT95), .B(new_n549), .C1(new_n551), .C2(new_n552), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G134gat), .B(G162gat), .Z(new_n561));
  NOR2_X1   g360(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n547), .B2(new_n549), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  OR2_X1    g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G57gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G64gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(G64gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(KEYINPUT88), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n574), .A2(new_n570), .A3(G64gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n569), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G64gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(G57gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT9), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n566), .A3(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G127gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n581), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n480), .B1(KEYINPUT21), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G155gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n590), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n547), .A2(new_n549), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n550), .A2(new_n555), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n563), .B(KEYINPUT90), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G120gat), .B(G148gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT99), .ZN(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n533), .A2(new_n581), .A3(new_n536), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n531), .A2(new_n588), .A3(new_n532), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n537), .A2(KEYINPUT10), .A3(new_n588), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n606), .B2(new_n608), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n605), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n612), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n609), .B2(new_n610), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT97), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n620), .B(new_n617), .C1(new_n609), .C2(new_n610), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n615), .A2(KEYINPUT98), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n605), .B1(new_n615), .B2(KEYINPUT98), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n616), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n565), .A2(new_n596), .A3(new_n600), .A4(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n514), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n256), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n470), .ZN(G1324gat));
  OAI21_X1  g430(.A(G8gat), .B1(new_n629), .B2(new_n319), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT100), .Z(new_n633));
  INV_X1    g432(.A(new_n629), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT16), .B(G8gat), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n318), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT42), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(G1325gat));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n373), .A2(KEYINPUT36), .ZN(new_n640));
  INV_X1    g439(.A(new_n426), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n425), .A2(KEYINPUT101), .A3(new_n426), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G15gat), .B1(new_n629), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n385), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n629), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n629), .A2(new_n343), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n625), .ZN(new_n652));
  INV_X1    g451(.A(new_n616), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n596), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n565), .A2(new_n600), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n514), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n453), .A3(new_n388), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n428), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n656), .A2(new_n509), .ZN(new_n666));
  INV_X1    g465(.A(new_n343), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n400), .B2(new_n421), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n644), .B1(new_n668), .B2(new_n389), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n658), .B1(new_n669), .B2(new_n387), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n665), .B(new_n666), .C1(new_n670), .C2(KEYINPUT44), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n643), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n425), .B2(new_n426), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n387), .B1(new_n423), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n657), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n663), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n679), .A2(KEYINPUT102), .A3(new_n665), .A4(new_n666), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n673), .A2(new_n388), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n662), .B1(new_n453), .B2(new_n681), .ZN(G1328gat));
  NAND3_X1  g481(.A1(new_n673), .A2(new_n680), .A3(new_n318), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G36gat), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n514), .A2(new_n449), .A3(new_n318), .A4(new_n659), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n690), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(G1329gat));
  AND3_X1   g491(.A1(new_n660), .A2(new_n459), .A3(new_n385), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n673), .A2(new_n680), .A3(new_n676), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G43gat), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n671), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n459), .B1(new_n699), .B2(new_n676), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n695), .A2(new_n696), .B1(new_n698), .B2(new_n700), .ZN(G1330gat));
  NAND2_X1  g500(.A1(new_n458), .A2(new_n460), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n660), .A2(new_n667), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n673), .A2(new_n680), .A3(new_n667), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n703), .B1(new_n699), .B2(new_n667), .ZN(new_n709));
  OAI22_X1  g508(.A1(KEYINPUT48), .A2(new_n706), .B1(new_n708), .B2(new_n709), .ZN(G1331gat));
  INV_X1    g509(.A(new_n596), .ZN(new_n711));
  NOR4_X1   g510(.A1(new_n657), .A2(new_n711), .A3(new_n508), .A4(new_n626), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n677), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n677), .A2(KEYINPUT105), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n256), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n570), .ZN(G1332gat));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n319), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  AND2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n723), .B(new_n726), .C1(new_n720), .C2(new_n721), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n717), .B2(new_n644), .ZN(new_n729));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n385), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n717), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1334gat));
  NOR2_X1   g533(.A1(new_n717), .A2(new_n343), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g535(.A1(new_n256), .A2(G85gat), .A3(new_n626), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n596), .A2(new_n508), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n678), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n670), .A2(KEYINPUT51), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n739), .A2(new_n654), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT107), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n679), .A2(new_n665), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n256), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n319), .A2(G92gat), .A3(new_n626), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G92gat), .B1(new_n749), .B2(new_n319), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n752), .B(KEYINPUT109), .Z(new_n756));
  NAND2_X1  g555(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(G1337gat));
  NOR3_X1   g559(.A1(new_n646), .A2(G99gat), .A3(new_n626), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT110), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n744), .B2(new_n745), .ZN(new_n763));
  OAI21_X1  g562(.A(G99gat), .B1(new_n749), .B2(new_n644), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1338gat));
  OAI21_X1  g564(.A(G106gat), .B1(new_n749), .B2(new_n343), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n343), .A2(G106gat), .A3(new_n626), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n743), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g569(.A1(new_n481), .A2(new_n483), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n496), .A2(new_n485), .A3(new_n497), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(new_n772), .B1(new_n441), .B2(new_n436), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n504), .A2(new_n505), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT86), .ZN(new_n775));
  INV_X1    g574(.A(new_n507), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n613), .A2(new_n620), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n609), .A2(new_n617), .A3(new_n610), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(KEYINPUT54), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n618), .A2(KEYINPUT97), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n783));
  AOI21_X1  g582(.A(new_n605), .B1(new_n618), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n784), .A3(KEYINPUT55), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n652), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n779), .A2(KEYINPUT54), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n619), .A2(new_n621), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n784), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND4_X1   g590(.A1(new_n657), .A2(new_n777), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n654), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n791), .A2(new_n508), .A3(new_n652), .A4(new_n785), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n657), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n711), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n565), .A2(new_n596), .A3(new_n600), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n798), .A2(new_n799), .A3(new_n509), .A4(new_n626), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT111), .B1(new_n627), .B2(new_n508), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n794), .A2(new_n793), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n658), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n657), .A2(new_n786), .A3(new_n777), .A4(new_n791), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n596), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n801), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT113), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n388), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n374), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n509), .A2(G113gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n319), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n667), .A2(new_n646), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n256), .A2(new_n318), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n809), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n513), .A3(new_n821), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n822), .A2(KEYINPUT115), .A3(G113gat), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT115), .B1(new_n822), .B2(G113gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n815), .B1(new_n823), .B2(new_n824), .ZN(G1340gat));
  NOR2_X1   g624(.A1(new_n626), .A2(G120gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n813), .A2(new_n319), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n654), .A3(new_n821), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(new_n829), .A3(G120gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(G120gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(G1341gat));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n319), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n596), .A2(new_n586), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n820), .A2(new_n596), .A3(new_n821), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n833), .A2(new_n834), .B1(new_n586), .B2(new_n835), .ZN(G1342gat));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n658), .A2(G134gat), .A3(new_n318), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n813), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n811), .A2(new_n812), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n810), .A2(KEYINPUT116), .A3(new_n374), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n820), .A2(new_n657), .A3(new_n821), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G134gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n843), .A3(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n809), .A2(new_n847), .A3(new_n667), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n782), .A2(new_n784), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n850));
  AOI22_X1  g649(.A1(new_n510), .A2(new_n512), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n851), .A2(new_n786), .B1(new_n654), .B2(new_n777), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n805), .B1(new_n852), .B2(new_n657), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n807), .B1(new_n853), .B2(new_n711), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT57), .B1(new_n854), .B2(new_n343), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n644), .A2(new_n817), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n848), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n508), .ZN(new_n859));
  INV_X1    g658(.A(new_n810), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n676), .A2(new_n343), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n318), .ZN(new_n863));
  INV_X1    g662(.A(new_n513), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(G141gat), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n859), .A2(G141gat), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n860), .A2(new_n319), .A3(new_n861), .A4(new_n865), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n867), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n205), .B1(new_n858), .B2(new_n513), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n866), .A2(new_n867), .B1(new_n869), .B2(new_n870), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n654), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n667), .A2(new_n847), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n711), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n864), .A2(new_n628), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n809), .A2(new_n667), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n872), .B(new_n876), .C1(new_n877), .C2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(G148gat), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT59), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n848), .A2(new_n855), .A3(new_n654), .A4(new_n856), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n203), .A2(KEYINPUT59), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT119), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n863), .A2(new_n203), .A3(new_n654), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1345gat));
  NOR3_X1   g686(.A1(new_n857), .A2(new_n208), .A3(new_n711), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n860), .A2(new_n319), .A3(new_n596), .A4(new_n861), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT120), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n890), .B2(new_n208), .ZN(G1346gat));
  OAI21_X1  g690(.A(G162gat), .B1(new_n857), .B2(new_n658), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n319), .A2(new_n657), .A3(new_n209), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n862), .B2(new_n893), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n319), .A2(new_n388), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n802), .A2(new_n808), .A3(new_n816), .A4(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT123), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(KEYINPUT123), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n513), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n802), .A2(new_n808), .A3(new_n256), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n802), .A2(new_n808), .A3(KEYINPUT121), .A4(new_n256), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n374), .A2(new_n319), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n908));
  INV_X1    g707(.A(new_n906), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n903), .B2(new_n904), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n509), .A2(new_n270), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n900), .A2(new_n261), .B1(new_n913), .B2(new_n914), .ZN(G1348gat));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n905), .B2(new_n906), .ZN(new_n917));
  AOI211_X1 g716(.A(KEYINPUT122), .B(new_n909), .C1(new_n903), .C2(new_n904), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n654), .A2(new_n262), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n654), .A3(new_n898), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G176gat), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n916), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT124), .B(new_n922), .C1(new_n913), .C2(new_n919), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n596), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G183gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n596), .A2(new_n280), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT125), .B1(new_n910), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n287), .B1(new_n899), .B2(new_n596), .ZN(new_n934));
  INV_X1    g733(.A(new_n932), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT60), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n897), .A2(new_n657), .A3(new_n898), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G190gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n941), .A3(G190gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n917), .A2(new_n918), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n658), .A2(G190gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT126), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947));
  INV_X1    g746(.A(new_n945), .ZN(new_n948));
  NOR4_X1   g747(.A1(new_n917), .A2(new_n918), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n943), .B1(new_n946), .B2(new_n949), .ZN(G1351gat));
  AOI21_X1  g749(.A(new_n876), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n644), .A3(new_n895), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(new_n864), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n676), .A2(new_n343), .A3(new_n319), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n905), .A2(new_n508), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n953), .B2(new_n956), .ZN(G1352gat));
  OAI21_X1  g756(.A(G204gat), .B1(new_n952), .B2(new_n626), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n626), .A2(G204gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n905), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(G1353gat));
  NAND4_X1  g762(.A1(new_n905), .A2(new_n302), .A3(new_n596), .A4(new_n955), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n644), .A2(new_n895), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n965), .B(new_n876), .C1(new_n877), .C2(KEYINPUT57), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n596), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  INV_X1    g768(.A(G211gat), .ZN(new_n970));
  AOI211_X1 g769(.A(new_n969), .B(new_n970), .C1(new_n966), .C2(new_n596), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n964), .B1(new_n968), .B2(new_n971), .ZN(G1354gat));
  AOI21_X1  g771(.A(new_n303), .B1(new_n966), .B2(new_n657), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n905), .A2(new_n303), .A3(new_n657), .A4(new_n955), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT127), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G218gat), .B1(new_n952), .B2(new_n658), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n978), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n979), .ZN(G1355gat));
endmodule


