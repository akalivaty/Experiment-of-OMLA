//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n582, new_n583, new_n584, new_n587, new_n589, new_n590, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  OAI211_X1 g037(.A(new_n462), .B(G125), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n467), .C1(new_n458), .C2(new_n459), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(G160));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(G136), .B2(new_n479), .ZN(G162));
  NOR2_X1   g055(.A1(new_n458), .A2(new_n459), .ZN(new_n481));
  NAND2_X1  g056(.A1(G126), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n481), .A2(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n458), .B2(new_n459), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n459), .C2(new_n458), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  XNOR2_X1  g069(.A(KEYINPUT6), .B(G651), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(G50), .A3(G543), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT67), .ZN(new_n497));
  INV_X1    g072(.A(G88), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT68), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n500), .A2(new_n503), .B1(KEYINPUT5), .B2(new_n499), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n495), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n497), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(G166));
  NAND2_X1  g085(.A1(new_n495), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G51), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n500), .A2(new_n503), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n518), .A2(new_n519), .A3(new_n495), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n517), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n508), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT69), .B(G90), .Z(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n505), .A2(new_n526), .B1(new_n527), .B2(new_n511), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  XNOR2_X1  g104(.A(KEYINPUT71), .B(G81), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n520), .A2(new_n530), .B1(new_n512), .B2(G43), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  NAND3_X1  g118(.A1(new_n495), .A2(G53), .A3(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT9), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT9), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n495), .A2(new_n546), .A3(G53), .A4(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n504), .A2(G91), .A3(new_n495), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n548), .B(new_n549), .C1(new_n508), .C2(new_n550), .ZN(G299));
  INV_X1    g126(.A(G171), .ZN(G301));
  INV_X1    g127(.A(G166), .ZN(G303));
  OAI21_X1  g128(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n512), .A2(G49), .ZN(new_n555));
  INV_X1    g130(.A(G87), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n505), .ZN(G288));
  NAND4_X1  g132(.A1(new_n518), .A2(G86), .A3(new_n519), .A4(new_n495), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n495), .A2(G48), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(G73), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n504), .B2(G61), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n558), .B(new_n559), .C1(new_n562), .C2(new_n508), .ZN(G305));
  AOI22_X1  g138(.A1(new_n520), .A2(G85), .B1(new_n512), .B2(G47), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT73), .Z(new_n565));
  AOI22_X1  g140(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n508), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G290));
  NAND2_X1  g143(.A1(G301), .A2(G868), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n520), .A2(G92), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT10), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G79), .A2(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(new_n519), .ZN(new_n574));
  INV_X1    g149(.A(G66), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n569), .B1(new_n579), .B2(G868), .ZN(G284));
  OAI21_X1  g155(.A(new_n569), .B1(new_n579), .B2(G868), .ZN(G321));
  NAND2_X1  g156(.A1(G286), .A2(G868), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT74), .Z(new_n583));
  INV_X1    g158(.A(G299), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(G868), .B2(new_n584), .ZN(G297));
  OAI21_X1  g160(.A(new_n583), .B1(G868), .B2(new_n584), .ZN(G280));
  INV_X1    g161(.A(G559), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n579), .B1(new_n587), .B2(G860), .ZN(G148));
  NAND2_X1  g163(.A1(new_n579), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G868), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g166(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g167(.A1(new_n467), .A2(G2104), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n471), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT13), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(G2100), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n479), .A2(G135), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n474), .A2(G123), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n467), .A2(G111), .ZN(new_n601));
  OAI21_X1  g176(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(G2096), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(G2096), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n598), .A2(new_n604), .A3(new_n605), .ZN(G156));
  XOR2_X1   g181(.A(G2451), .B(G2454), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT16), .ZN(new_n608));
  XNOR2_X1  g183(.A(G1341), .B(G1348), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT75), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT14), .ZN(new_n612));
  XNOR2_X1  g187(.A(G2427), .B(G2438), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2430), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT15), .B(G2435), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(new_n614), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n611), .B(new_n617), .Z(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2443), .B(G2446), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(G14), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n619), .ZN(G401));
  XOR2_X1   g198(.A(G2084), .B(G2090), .Z(new_n624));
  XNOR2_X1  g199(.A(G2067), .B(G2678), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2072), .B(G2078), .Z(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT77), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT76), .B(KEYINPUT18), .Z(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  OAI21_X1  g207(.A(KEYINPUT17), .B1(new_n624), .B2(new_n625), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(new_n627), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n627), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(new_n626), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2096), .B(G2100), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(G227));
  XNOR2_X1  g214(.A(G1971), .B(G1976), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT19), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1961), .B(G1966), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT78), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1956), .B(G2474), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n646), .A3(new_n641), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n647), .B1(new_n646), .B2(new_n641), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1991), .B(G1996), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1981), .B(G1986), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(G229));
  NAND2_X1  g235(.A1(new_n474), .A2(G129), .ZN(new_n661));
  NAND3_X1  g236(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT26), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n664), .A2(new_n665), .B1(G105), .B2(new_n594), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(G141), .B2(new_n479), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G29), .ZN(new_n669));
  NOR2_X1   g244(.A1(G29), .A2(G32), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(KEYINPUT92), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(KEYINPUT92), .B2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT27), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n467), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT91), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n479), .A2(G139), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT90), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(G33), .B(new_n683), .S(G29), .Z(new_n684));
  AND2_X1   g259(.A1(new_n684), .A2(G2072), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(G2072), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT80), .B(G29), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(G27), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G164), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  INV_X1    g266(.A(G2078), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NOR2_X1   g269(.A1(G171), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G5), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR4_X1   g273(.A1(new_n685), .A2(new_n686), .A3(new_n693), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n674), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G168), .A2(new_n694), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n694), .B2(G21), .ZN(new_n702));
  INV_X1    g277(.A(G1966), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT31), .B(G11), .Z(new_n706));
  INV_X1    g281(.A(G28), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT93), .Z(new_n709));
  AOI21_X1  g284(.A(G29), .B1(new_n707), .B2(KEYINPUT30), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n603), .B2(new_n687), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n703), .B2(new_n702), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT24), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G34), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(G34), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n688), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G160), .B2(G29), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n696), .A2(new_n697), .B1(G2084), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n691), .A2(new_n692), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n720), .B(new_n721), .C1(G2084), .C2(new_n719), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n700), .A2(new_n714), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n687), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n474), .A2(G128), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT86), .Z(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G116), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n479), .A2(G140), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n727), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT88), .B(G2067), .Z(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n579), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G4), .B2(G16), .ZN(new_n744));
  INV_X1    g319(.A(G1348), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n740), .A2(new_n741), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n742), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n688), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n688), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2090), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n694), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT23), .Z(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1956), .Z(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G19), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n537), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1341), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n749), .A2(new_n753), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n725), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G22), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G166), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G1971), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(G16), .A2(G23), .ZN(new_n767));
  OR2_X1    g342(.A1(G288), .A2(KEYINPUT84), .ZN(new_n768));
  NAND2_X1  g343(.A1(G288), .A2(KEYINPUT84), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n767), .B1(new_n770), .B2(new_n694), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT33), .B(G1976), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n694), .A2(G6), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n518), .A2(G61), .A3(new_n519), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n508), .B1(new_n776), .B2(new_n560), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n558), .A2(new_n559), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n775), .B1(new_n779), .B2(new_n694), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n766), .A2(new_n773), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n479), .A2(G131), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n474), .A2(G119), .ZN(new_n786));
  OR2_X1    g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G25), .B(new_n789), .S(new_n688), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT82), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT35), .B(G1991), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT81), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G24), .ZN(new_n796));
  INV_X1    g371(.A(G290), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT83), .B(G1986), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n784), .A2(new_n794), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT85), .B(KEYINPUT36), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n724), .B(new_n762), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT85), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n803), .A2(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  NAND2_X1  g383(.A1(new_n579), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n508), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n505), .A2(new_n813), .B1(new_n814), .B2(new_n511), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n536), .B(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n810), .B(new_n817), .Z(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n819));
  INV_X1    g394(.A(G860), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  INV_X1    g400(.A(new_n482), .ZN(new_n826));
  INV_X1    g401(.A(new_n486), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n471), .A2(new_n826), .B1(new_n827), .B2(new_n484), .ZN(new_n828));
  INV_X1    g403(.A(new_n493), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n492), .B1(new_n471), .B2(new_n489), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n491), .A2(new_n493), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(KEYINPUT96), .A3(new_n828), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n737), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n479), .A2(G142), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n474), .A2(G130), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n467), .A2(G118), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n789), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n596), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n668), .B(new_n683), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n603), .B(G160), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(G162), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT98), .B(G37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g430(.A(new_n589), .B(new_n817), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n578), .A2(new_n584), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n579), .A2(G299), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n857), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(KEYINPUT41), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n865), .B2(new_n856), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(G290), .B(new_n770), .ZN(new_n871));
  XNOR2_X1  g446(.A(G166), .B(G305), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n873), .A3(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G868), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n879));
  INV_X1    g454(.A(new_n816), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(G868), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G868), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n875), .B2(new_n876), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT100), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(G295));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n882), .ZN(G331));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n817), .B(G301), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(G168), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(G168), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n865), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(new_n861), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n889), .B1(new_n898), .B2(new_n874), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n873), .B1(new_n894), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(KEYINPUT41), .A3(new_n864), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n873), .B(new_n902), .C1(new_n903), .C2(new_n861), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n874), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n853), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(KEYINPUT43), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n899), .B2(new_n900), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n908), .B2(new_n906), .ZN(new_n910));
  MUX2_X1   g485(.A(new_n907), .B(new_n910), .S(KEYINPUT44), .Z(G397));
  INV_X1    g486(.A(KEYINPUT126), .ZN(new_n912));
  INV_X1    g487(.A(G1384), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n836), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n469), .A2(G40), .A3(new_n468), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n466), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1996), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT46), .ZN(new_n923));
  INV_X1    g498(.A(G2067), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n737), .B(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(new_n668), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n920), .B(KEYINPUT102), .Z(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n923), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT47), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n925), .B1(new_n921), .B2(new_n668), .ZN(new_n931));
  INV_X1    g506(.A(new_n922), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n931), .A2(new_n927), .B1(new_n668), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n792), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n789), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n789), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n927), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1986), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n797), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT101), .Z(new_n941));
  INV_X1    g516(.A(new_n920), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT48), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n930), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n933), .A2(new_n936), .B1(new_n924), .B2(new_n738), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n928), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT63), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT45), .B1(new_n831), .B2(new_n913), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n919), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n915), .A2(G1384), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n833), .A2(new_n835), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G1971), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G2090), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n917), .B1(new_n465), .B2(G2105), .ZN(new_n957));
  XOR2_X1   g532(.A(KEYINPUT103), .B(KEYINPUT50), .Z(new_n958));
  AOI211_X1 g533(.A(G1384), .B(new_n958), .C1(new_n834), .C2(new_n828), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT50), .B1(new_n831), .B2(new_n913), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n956), .B(new_n957), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n950), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(G166), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT55), .B(G8), .C1(new_n506), .C2(new_n509), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n833), .A2(new_n835), .A3(new_n953), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n834), .B2(new_n828), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n957), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n765), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT104), .A3(new_n961), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n963), .A2(G8), .A3(new_n968), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT105), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n831), .A2(new_n913), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n915), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n954), .A2(new_n957), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(G164), .B2(G1384), .ZN(new_n980));
  INV_X1    g555(.A(new_n958), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n831), .A2(new_n913), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n919), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n978), .A2(new_n765), .B1(new_n983), .B2(new_n956), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n965), .B1(new_n984), .B2(KEYINPUT104), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n968), .A4(new_n963), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n768), .A2(G1976), .A3(new_n769), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n965), .B1(new_n957), .B2(new_n970), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT52), .ZN(new_n992));
  INV_X1    g567(.A(G1976), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(G288), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(G305), .B2(G1981), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n998));
  INV_X1    g573(.A(G1981), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n779), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n778), .A2(KEYINPUT107), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n558), .A2(new_n1002), .A3(new_n559), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1001), .B(new_n1003), .C1(new_n508), .C2(new_n562), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n997), .A2(new_n1000), .B1(new_n1004), .B2(G1981), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n990), .B1(new_n1005), .B2(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n997), .A2(new_n1000), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(G1981), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT108), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n990), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n996), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n968), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n831), .A2(new_n979), .A3(new_n913), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n957), .C1(new_n970), .C2(new_n958), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2090), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n955), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n988), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1025));
  AOI211_X1 g600(.A(G2084), .B(new_n917), .C1(new_n465), .C2(G2105), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n959), .B2(new_n960), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n831), .A2(new_n953), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n957), .C1(new_n970), .C2(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n703), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT111), .B(new_n1026), .C1(new_n959), .C2(new_n960), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(G8), .A3(G168), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n949), .B1(new_n1025), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n968), .B1(new_n985), .B2(new_n963), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1037), .A2(new_n1035), .A3(new_n949), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(new_n1018), .A3(new_n988), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1018), .A2(new_n975), .A3(new_n987), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n990), .B(KEYINPUT109), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G288), .A2(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1015), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1006), .A2(new_n1009), .A3(KEYINPUT108), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1007), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(KEYINPUT110), .A3(new_n1007), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1041), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G78), .A2(G543), .ZN(new_n1052));
  INV_X1    g627(.A(G65), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n574), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1054), .A2(G651), .B1(G91), .B2(new_n520), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n548), .C1(KEYINPUT113), .C2(KEYINPUT57), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT113), .B(new_n549), .C1(new_n550), .C2(new_n508), .ZN(new_n1058));
  NAND3_X1  g633(.A1(G299), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT112), .B(G1956), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1021), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n954), .A2(new_n977), .A3(new_n957), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n980), .A2(new_n982), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n957), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n745), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n957), .A2(new_n970), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(new_n957), .B2(new_n970), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n924), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n578), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1060), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1065), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1065), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1060), .A2(new_n1062), .A3(KEYINPUT117), .A4(new_n1064), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT61), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1078), .A2(KEYINPUT118), .A3(KEYINPUT61), .A4(new_n1079), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AND4_X1   g659(.A1(KEYINPUT60), .A2(new_n1068), .A3(new_n1073), .A4(new_n578), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n919), .B2(new_n976), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1070), .A3(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n954), .A2(new_n977), .A3(new_n921), .A4(new_n957), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT59), .B1(new_n1090), .B2(new_n537), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1092), .B(new_n536), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1085), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1068), .A2(new_n1073), .A3(KEYINPUT60), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n579), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1060), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1065), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT115), .B(KEYINPUT61), .Z(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT116), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1104), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1106), .B(new_n1107), .C1(new_n1102), .C2(new_n1065), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1094), .B(new_n1099), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1076), .B1(new_n1084), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT111), .B1(new_n1066), .B2(new_n1026), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1029), .A2(KEYINPUT119), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(G168), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n965), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G286), .A2(G8), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1034), .B2(G8), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1120), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(KEYINPUT120), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1122), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n978), .B2(G2078), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1067), .A2(new_n697), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n692), .A2(KEYINPUT53), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n916), .A2(new_n957), .A3(new_n1136), .A4(new_n954), .ZN(new_n1137));
  AOI21_X1  g712(.A(G301), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n952), .A2(new_n1030), .A3(new_n1136), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1133), .A2(new_n1139), .A3(new_n1134), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n1140), .B2(G171), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(G171), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1135), .A2(G301), .A3(new_n1137), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1110), .A2(new_n1131), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1025), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n975), .A2(new_n987), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(KEYINPUT123), .A3(new_n1018), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1040), .B(new_n1051), .C1(new_n1150), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1127), .A2(new_n1157), .A3(new_n1130), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1152), .A3(new_n1159), .A4(new_n1154), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT120), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1129), .A2(new_n1128), .A3(new_n1125), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT62), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT125), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1131), .A2(new_n1166), .A3(KEYINPUT62), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1156), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n941), .B1(new_n939), .B2(new_n797), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n920), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n937), .A3(new_n933), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n912), .B(new_n948), .C1(new_n1171), .C2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1025), .A2(new_n1151), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT123), .B1(new_n1153), .B2(new_n1018), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1166), .B1(new_n1131), .B2(KEYINPUT62), .ZN(new_n1181));
  AOI211_X1 g756(.A(KEYINPUT125), .B(new_n1157), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1180), .A2(new_n1183), .A3(new_n1170), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1051), .A2(new_n1040), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1174), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n945), .A2(new_n947), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT126), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1175), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g766(.A(G229), .ZN(new_n1193));
  INV_X1    g767(.A(G319), .ZN(new_n1194));
  NOR3_X1   g768(.A1(G401), .A2(new_n1194), .A3(G227), .ZN(new_n1195));
  XOR2_X1   g769(.A(new_n1195), .B(KEYINPUT127), .Z(new_n1196));
  NAND4_X1  g770(.A1(new_n907), .A2(new_n1193), .A3(new_n854), .A4(new_n1196), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


