//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT64), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G50), .B(G68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XOR2_X1   g0034(.A(G58), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  NAND2_X1  g0040(.A1(G33), .A2(G41), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n241), .A2(G1), .A3(G13), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G274), .ZN(new_n243));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n242), .ZN(new_n247));
  INV_X1    g0047(.A(new_n245), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n246), .B1(G226), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(G223), .B1(new_n259), .B2(G77), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1698), .B1(new_n254), .B2(new_n255), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G222), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n250), .B1(new_n263), .B2(new_n242), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G169), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n211), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n212), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n212), .B1(new_n201), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n273), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G50), .ZN(new_n287));
  INV_X1    g0087(.A(new_n273), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n244), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n287), .B1(new_n291), .B2(G50), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n284), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n268), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n271), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n269), .A2(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n268), .A2(G190), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n293), .B(KEYINPUT9), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n298), .A2(new_n303), .A3(new_n299), .A4(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n297), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G97), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n253), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n261), .B2(G226), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n254), .A2(new_n255), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G232), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n251), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n247), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n246), .B1(G238), .B2(new_n249), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G190), .ZN(new_n319));
  INV_X1    g0119(.A(new_n317), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G200), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT71), .B1(new_n286), .B2(G68), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n288), .A2(G68), .A3(new_n286), .A4(new_n289), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n278), .A2(new_n280), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n275), .A2(new_n327), .B1(new_n212), .B2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n273), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n325), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n324), .B(new_n331), .C1(new_n330), .C2(new_n329), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n319), .A2(new_n322), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n332), .B(KEYINPUT72), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT14), .B1(new_n318), .B2(new_n270), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n318), .A2(G179), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n321), .A2(new_n338), .A3(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n334), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT15), .B(G87), .Z(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n275), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n274), .A2(new_n278), .B1(new_n212), .B2(new_n327), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n273), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n291), .A2(G77), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n346), .B(new_n347), .C1(G77), .C2(new_n286), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n256), .A2(G238), .B1(new_n259), .B2(G107), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(G1698), .B2(new_n310), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n247), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n246), .B1(G244), .B2(new_n249), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(KEYINPUT68), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT68), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n348), .B1(new_n357), .B2(G200), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n353), .B(KEYINPUT68), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT69), .B1(new_n359), .B2(G190), .ZN(new_n360));
  OAI211_X1 g0160(.A(KEYINPUT69), .B(G190), .C1(new_n354), .C2(new_n356), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n294), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n357), .A2(new_n270), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n348), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n305), .B(new_n341), .C1(new_n367), .C2(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT70), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  AND2_X1   g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT73), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(G20), .C1(new_n371), .C2(new_n201), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n277), .A2(G159), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G68), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n309), .B2(G20), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n370), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n259), .B2(new_n212), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n257), .A2(new_n258), .A3(new_n380), .A4(G20), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n373), .A2(new_n375), .B1(G159), .B2(new_n277), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n273), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n274), .ZN(new_n391));
  INV_X1    g0191(.A(new_n286), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n391), .B2(new_n290), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(G223), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n397));
  OAI211_X1 g0197(.A(G226), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n398));
  INV_X1    g0198(.A(G87), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n397), .B(new_n398), .C1(new_n253), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n247), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n242), .A2(G232), .A3(new_n245), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n243), .B2(new_n245), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G169), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n400), .B2(new_n247), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n396), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n390), .A2(new_n395), .B1(new_n406), .B2(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G190), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(new_n415), .A3(new_n404), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G200), .B2(new_n407), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n390), .A2(new_n417), .A3(new_n395), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n387), .A2(new_n388), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n288), .B1(new_n421), .B2(new_n370), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n394), .B1(new_n422), .B2(new_n389), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n417), .ZN(new_n424));
  AND4_X1   g0224(.A1(new_n411), .A2(new_n414), .A3(new_n420), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n369), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n368), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n286), .A2(G116), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n244), .A2(G33), .ZN(new_n429));
  AND4_X1   g0229(.A1(new_n211), .A2(new_n286), .A3(new_n272), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(G116), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n432));
  OAI21_X1  g0232(.A(new_n212), .B1(new_n306), .B2(G33), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(G33), .A3(G283), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G283), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT75), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n273), .B1(new_n212), .B2(G116), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G116), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n272), .A2(new_n211), .B1(G20), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n437), .A2(new_n435), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n433), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n431), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT21), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  INV_X1    g0250(.A(new_n211), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n448), .A2(new_n450), .B1(new_n451), .B2(new_n241), .ZN(new_n452));
  INV_X1    g0252(.A(G274), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n451), .B2(new_n241), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n244), .A2(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n452), .A2(G270), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G257), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n461));
  OAI211_X1 g0261(.A(G264), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n254), .A2(G303), .A3(new_n255), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n247), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n447), .B(new_n270), .C1(new_n460), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n465), .A3(G179), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n446), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n460), .A2(new_n465), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n446), .B1(G200), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n415), .B2(new_n470), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n446), .A3(G169), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT84), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n473), .A2(new_n474), .A3(new_n447), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n473), .B2(new_n447), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n469), .B(new_n472), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT85), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n447), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n474), .A3(new_n447), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(KEYINPUT85), .A3(new_n469), .A4(new_n472), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n253), .A2(new_n441), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n261), .B2(G238), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT77), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n256), .B2(G244), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(KEYINPUT77), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT78), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n256), .A2(new_n488), .A3(G244), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(KEYINPUT77), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT78), .A3(new_n487), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n242), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n455), .A2(G250), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n454), .A2(new_n450), .B1(new_n500), .B2(new_n242), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G200), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n497), .A2(KEYINPUT78), .A3(new_n487), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT78), .B1(new_n497), .B2(new_n487), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n247), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G190), .A3(new_n501), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n342), .A2(new_n286), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n275), .B2(new_n306), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n309), .A2(new_n212), .A3(G68), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT79), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G87), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n523));
  XNOR2_X1  g0323(.A(KEYINPUT79), .B(G87), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(new_n521), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(new_n307), .B2(KEYINPUT19), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n517), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI211_X1 g0330(.A(KEYINPUT81), .B(new_n528), .C1(new_n523), .C2(new_n526), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n516), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n508), .B1(new_n532), .B2(new_n273), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n288), .A2(new_n286), .A3(new_n429), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n430), .A2(KEYINPUT74), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G87), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n503), .A2(new_n507), .A3(new_n533), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n508), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n342), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n527), .A2(new_n529), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT81), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n527), .A2(new_n517), .A3(new_n529), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n515), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n541), .B(new_n542), .C1(new_n546), .C2(new_n288), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n270), .B1(new_n499), .B2(new_n502), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n506), .A2(new_n294), .A3(new_n501), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n540), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n486), .A2(new_n212), .ZN(new_n552));
  INV_X1    g0352(.A(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT23), .B1(new_n553), .B2(G20), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT23), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n555), .A2(new_n212), .A3(G107), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n212), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT22), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n309), .A2(new_n560), .A3(new_n212), .A4(G87), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g0362(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n563), .B(new_n557), .C1(new_n559), .C2(new_n561), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n273), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n392), .A2(KEYINPUT25), .A3(new_n553), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT87), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT25), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n286), .B2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT88), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n538), .A2(G107), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n309), .A2(G257), .A3(G1698), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  OAI211_X1 g0376(.A(G250), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n247), .B1(G264), .B2(new_n452), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n459), .A2(new_n454), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n270), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(KEYINPUT89), .B1(new_n582), .B2(new_n294), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(KEYINPUT89), .A3(G169), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n574), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n582), .A2(G190), .ZN(new_n586));
  AOI21_X1  g0386(.A(G200), .B1(new_n579), .B2(new_n580), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n567), .B(new_n573), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  AND2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n521), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n553), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n594), .A2(new_n212), .B1(new_n327), .B2(new_n278), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n553), .B1(new_n381), .B2(new_n382), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n273), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n536), .A2(new_n537), .A3(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n392), .A2(new_n306), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n458), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n450), .B1(new_n601), .B2(new_n456), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G257), .A3(new_n242), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n580), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G244), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT4), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n309), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n437), .A2(new_n435), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n309), .A2(G250), .A3(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n611), .B2(new_n247), .ZN(new_n612));
  INV_X1    g0412(.A(G200), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n600), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n247), .ZN(new_n616));
  INV_X1    g0416(.A(new_n604), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT76), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT76), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(G190), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  AOI211_X1 g0423(.A(KEYINPUT76), .B(new_n604), .C1(new_n247), .C2(new_n611), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n616), .B2(new_n617), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n270), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G107), .B1(new_n385), .B2(new_n386), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n592), .A2(new_n593), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n630), .A2(new_n273), .B1(new_n306), .B2(new_n392), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n598), .B1(new_n294), .B2(new_n612), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n551), .A2(new_n589), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n427), .A2(new_n485), .A3(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n506), .A2(KEYINPUT90), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n499), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n502), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n549), .B(new_n547), .C1(new_n640), .C2(G169), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n626), .A2(new_n632), .A3(KEYINPUT91), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT91), .B1(new_n626), .B2(new_n632), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n533), .A2(new_n539), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n507), .B(new_n645), .C1(new_n640), .C2(new_n613), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n641), .A2(new_n644), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n585), .A2(new_n469), .A3(new_n483), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n623), .A2(new_n633), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n646), .A2(new_n649), .A3(new_n650), .A4(new_n588), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT26), .B1(new_n551), .B2(new_n633), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n648), .A2(new_n641), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n427), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n412), .B(KEYINPUT18), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n340), .A2(new_n335), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n366), .B2(new_n334), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n420), .A2(new_n424), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n302), .A2(new_n304), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n297), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n654), .A2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n244), .A2(new_n212), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n446), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n479), .B2(new_n484), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n483), .A2(new_n469), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n672), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n670), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n567), .B2(new_n573), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n589), .A2(new_n681), .B1(new_n585), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n585), .A2(new_n670), .ZN(new_n684));
  INV_X1    g0484(.A(new_n589), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n670), .B1(new_n483), .B2(new_n469), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n527), .A2(G116), .ZN(new_n689));
  INV_X1    g0489(.A(new_n206), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n209), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n653), .A2(new_n680), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n647), .ZN(new_n701));
  INV_X1    g0501(.A(new_n633), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n540), .A3(new_n550), .A4(new_n647), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n651), .A2(new_n703), .A3(new_n641), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT29), .B(new_n680), .C1(new_n701), .C2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n701), .A2(new_n704), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT94), .A3(KEYINPUT29), .A4(new_n680), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n670), .B1(new_n479), .B2(new_n484), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n635), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n578), .A2(new_n247), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n452), .A2(G264), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n467), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n506), .A2(new_n716), .A3(new_n501), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n619), .A2(new_n621), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n499), .A2(new_n502), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n624), .A2(new_n625), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT30), .A4(new_n716), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n460), .B2(new_n465), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n618), .A2(new_n582), .A3(KEYINPUT93), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT93), .B1(new_n618), .B2(new_n582), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n719), .B(new_n722), .C1(new_n640), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n670), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g0530(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n731));
  OAI211_X1 g0531(.A(new_n711), .B(new_n730), .C1(new_n728), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n709), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n695), .B1(new_n735), .B2(G1), .ZN(G364));
  AND2_X1   g0536(.A1(new_n212), .A2(G13), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n244), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n691), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n679), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n677), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(G330), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT98), .Z(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n677), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n740), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n212), .A2(new_n294), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n415), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n753), .A2(G68), .B1(new_n754), .B2(G50), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G20), .A3(new_n294), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G159), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT32), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n212), .A2(new_n613), .A3(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n755), .B(new_n760), .C1(new_n524), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n415), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n415), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n212), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(G107), .B1(new_n768), .B2(G97), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(KEYINPUT32), .B2(new_n759), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n751), .A2(new_n756), .ZN(new_n771));
  INV_X1    g0571(.A(G58), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n751), .A2(G190), .A3(new_n613), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n309), .B1(new_n771), .B2(new_n327), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n763), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n773), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G322), .B1(G329), .B2(new_n758), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n259), .C1(new_n778), .C2(new_n771), .ZN(new_n779));
  INV_X1    g0579(.A(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n753), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n754), .A2(G326), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n762), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n764), .A2(new_n787), .B1(new_n767), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n779), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n775), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n211), .B1(G20), .B2(new_n270), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n750), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n748), .A2(new_n792), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n309), .A2(new_n206), .ZN(new_n796));
  INV_X1    g0596(.A(G355), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n797), .B1(G116), .B2(new_n206), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT95), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n259), .A2(new_n206), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT96), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n449), .B2(new_n210), .ZN(new_n803));
  INV_X1    g0603(.A(new_n236), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(KEYINPUT97), .B1(new_n804), .B2(G45), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n799), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n749), .B(new_n793), .C1(new_n795), .C2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n743), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  INV_X1    g0610(.A(new_n366), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n680), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT69), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n357), .B2(new_n415), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n361), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(new_n358), .B1(new_n348), .B2(new_n670), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n812), .B1(new_n816), .B2(new_n811), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n696), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n366), .A2(new_n670), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n348), .A2(new_n670), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n363), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n821), .B2(new_n366), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n653), .A2(new_n822), .A3(new_n680), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n740), .B1(new_n824), .B2(new_n733), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n733), .B2(new_n824), .ZN(new_n826));
  INV_X1    g0626(.A(new_n771), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n776), .A2(G143), .B1(new_n827), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(new_n754), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(new_n753), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n828), .B1(new_n829), .B2(new_n830), .C1(new_n276), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n765), .A2(G68), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n309), .C1(new_n837), .C2(new_n757), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n762), .A2(new_n280), .B1(new_n767), .B2(new_n772), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n834), .A2(new_n835), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n829), .A2(new_n785), .B1(new_n553), .B2(new_n762), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G97), .A2(new_n768), .B1(new_n753), .B2(G283), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n309), .B1(new_n776), .B2(G294), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n827), .A2(G116), .B1(new_n758), .B2(G311), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n841), .B(new_n845), .C1(G87), .C2(new_n765), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n792), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n792), .A2(new_n744), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n750), .B1(new_n327), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n822), .C2(new_n745), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n826), .A2(new_n850), .ZN(G384));
  NAND2_X1  g0651(.A1(new_n335), .A2(new_n670), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n657), .A2(new_n333), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n335), .B(new_n670), .C1(new_n334), .C2(new_n340), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(new_n822), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT105), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n858));
  INV_X1    g0658(.A(new_n731), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n727), .B2(new_n670), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n861), .B2(new_n711), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n728), .A2(new_n731), .ZN(new_n864));
  AND4_X1   g0664(.A1(new_n857), .A2(new_n711), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n856), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n668), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n396), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n655), .B2(new_n659), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT101), .ZN(new_n872));
  INV_X1    g0672(.A(new_n409), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n418), .B1(new_n423), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n423), .B2(new_n668), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n872), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT37), .B1(new_n396), .B2(new_n869), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(KEYINPUT101), .A3(new_n410), .A4(new_n418), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n410), .A2(new_n870), .A3(new_n418), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n877), .A2(new_n879), .B1(KEYINPUT37), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n871), .B1(new_n881), .B2(KEYINPUT103), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n879), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n868), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT16), .B1(new_n387), .B2(new_n388), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT99), .B1(new_n889), .B2(new_n288), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT99), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n384), .A2(new_n891), .A3(new_n273), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n892), .A3(new_n389), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n395), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT100), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n896), .A3(new_n395), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n869), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT38), .B1(new_n425), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n895), .A2(new_n409), .A3(new_n897), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n900), .A3(new_n418), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(new_n883), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT40), .B1(new_n888), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT106), .B1(new_n866), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  INV_X1    g0706(.A(new_n871), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n885), .B2(new_n886), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n867), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n899), .ZN(new_n911));
  INV_X1    g0711(.A(new_n418), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n893), .A2(new_n896), .A3(new_n395), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n896), .B1(new_n893), .B2(new_n395), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n915), .B2(new_n409), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n875), .B1(new_n916), .B2(new_n898), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n877), .A2(new_n879), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n906), .B1(new_n910), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n855), .A2(new_n822), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n864), .A2(new_n863), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n635), .A2(new_n710), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT105), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n861), .A2(new_n857), .A3(new_n711), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n920), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n918), .B1(new_n901), .B2(KEYINPUT37), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n425), .A2(new_n898), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n919), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n905), .A2(new_n928), .B1(new_n906), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n426), .B(new_n368), .C1(new_n925), .C2(new_n924), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n678), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n340), .A2(new_n335), .A3(new_n680), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n910), .A2(new_n919), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n932), .B2(new_n919), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n855), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n823), .B2(new_n812), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n948), .A2(new_n933), .B1(new_n656), .B2(new_n668), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n706), .A2(new_n708), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n427), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n663), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n951), .B(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n939), .A2(new_n955), .B1(new_n244), .B2(new_n737), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n939), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n628), .A2(KEYINPUT35), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n628), .A2(KEYINPUT35), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n958), .A2(G116), .A3(new_n213), .A4(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT36), .Z(new_n961));
  OR3_X1    g0761(.A1(new_n209), .A2(new_n327), .A3(new_n371), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n280), .A2(G68), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n244), .B(G13), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n957), .A2(new_n961), .A3(new_n964), .ZN(G367));
  INV_X1    g0765(.A(new_n683), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n600), .A2(new_n670), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n650), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n702), .A2(new_n670), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT107), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n684), .A4(new_n687), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n687), .A2(new_n684), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT107), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n971), .A2(new_n975), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT44), .Z(new_n981));
  NAND3_X1  g0781(.A1(new_n974), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n967), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n687), .B1(new_n682), .B2(new_n686), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n679), .B(new_n987), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n709), .A2(new_n733), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT108), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n985), .A2(new_n986), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n734), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n691), .B(KEYINPUT41), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n738), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n971), .A2(new_n687), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  INV_X1    g0798(.A(new_n623), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n633), .B1(new_n999), .B2(new_n585), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n997), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n645), .A2(new_n680), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n641), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n641), .A2(new_n646), .A3(new_n1002), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n998), .A2(new_n1001), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n966), .A2(new_n972), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n996), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1003), .A2(new_n748), .A3(new_n1004), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n794), .B1(new_n206), .B2(new_n343), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n231), .B2(new_n801), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n765), .A2(G77), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n309), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT110), .Z(new_n1017));
  OAI22_X1  g0817(.A1(new_n773), .A2(new_n276), .B1(new_n771), .B2(new_n280), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G137), .B2(new_n758), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G68), .A2(new_n768), .B1(new_n753), .B2(G159), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n762), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G58), .A2(new_n1021), .B1(new_n754), .B2(G143), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G107), .A2(new_n768), .B1(new_n754), .B2(G311), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n306), .B2(new_n764), .C1(new_n788), .C2(new_n831), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n776), .A2(G303), .B1(G317), .B2(new_n758), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT46), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n762), .B2(new_n441), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n309), .B1(new_n827), .B2(G283), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1017), .A2(new_n1023), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n750), .B(new_n1014), .C1(new_n1033), .C2(new_n792), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1012), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1011), .A2(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n734), .A2(new_n988), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1037), .A2(new_n691), .A3(new_n990), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n228), .A2(G45), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n274), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g0841(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n689), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n801), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n689), .A2(new_n796), .B1(G107), .B2(new_n206), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT111), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1044), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n740), .B1(new_n1049), .B2(new_n795), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n682), .A2(new_n747), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n827), .A2(G68), .B1(new_n758), .B2(G150), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n309), .C1(new_n280), .C2(new_n773), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1021), .A2(G77), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n768), .A2(new_n342), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n274), .C2(new_n831), .ZN(new_n1056));
  INV_X1    g0856(.A(G159), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n829), .A2(new_n1057), .B1(new_n306), .B2(new_n764), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1053), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT112), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n309), .B1(new_n758), .B2(G326), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n762), .A2(new_n788), .B1(new_n767), .B2(new_n787), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n776), .A2(G317), .B1(new_n827), .B2(G303), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n754), .A2(G322), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n778), .C2(new_n831), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1061), .B1(new_n441), .B2(new_n764), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1060), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1050), .B(new_n1051), .C1(new_n792), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n989), .B2(new_n739), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1038), .A2(new_n1074), .ZN(G393));
  XOR2_X1   g0875(.A(new_n983), .B(new_n984), .Z(new_n1076));
  AOI21_X1  g0876(.A(new_n692), .B1(new_n1076), .B2(new_n990), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n992), .A2(new_n993), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1076), .A2(new_n738), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n829), .A2(new_n276), .B1(new_n1057), .B2(new_n773), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n767), .A2(new_n327), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n259), .B1(new_n758), .B2(G143), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n399), .B2(new_n764), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(G68), .C2(new_n1021), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n753), .A2(G50), .B1(new_n827), .B2(new_n391), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT113), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1082), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G317), .A2(new_n754), .B1(new_n776), .B2(G311), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n831), .A2(new_n785), .B1(new_n553), .B2(new_n764), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n309), .B1(new_n758), .B2(G322), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n788), .B2(new_n771), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n762), .A2(new_n787), .B1(new_n767), .B2(new_n441), .ZN(new_n1097));
  OR3_X1    g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1091), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n792), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n795), .B1(G97), .B2(new_n690), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n801), .A2(new_n239), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n750), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n972), .C2(new_n747), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1079), .A2(new_n1080), .A3(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n933), .A2(KEYINPUT39), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n910), .A2(new_n919), .A3(new_n942), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n941), .C2(new_n948), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n821), .A2(new_n366), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n680), .B(new_n1110), .C1(new_n701), .C2(new_n704), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n812), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n855), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n941), .B1(new_n910), .B2(new_n919), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n856), .C1(new_n862), .C2(new_n865), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT115), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n678), .B1(new_n924), .B2(new_n925), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT115), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n856), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n732), .A2(G330), .A3(new_n822), .A4(new_n855), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1126), .A2(new_n1109), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1126), .B2(new_n1109), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1123), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1125), .A2(new_n1112), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n678), .B(new_n817), .C1(new_n924), .C2(new_n925), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(KEYINPUT117), .C1(new_n855), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n855), .B1(new_n1119), .B2(new_n822), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1124), .A2(new_n812), .A3(new_n1111), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n947), .B1(new_n733), .B2(new_n817), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1118), .A2(new_n1121), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n823), .A2(new_n812), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n427), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n953), .A2(new_n663), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1131), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n692), .B1(new_n1149), .B2(new_n1130), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1131), .A2(new_n739), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1107), .A2(new_n744), .A3(new_n1108), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n553), .A2(new_n831), .B1(new_n829), .B2(new_n787), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G87), .B2(new_n1021), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1083), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n773), .A2(new_n441), .B1(new_n771), .B2(new_n306), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n309), .B(new_n1157), .C1(G294), .C2(new_n758), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n836), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1021), .A2(G150), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT118), .Z(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n827), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n309), .B1(new_n773), .B2(new_n837), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G125), .B2(new_n758), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G159), .A2(new_n768), .B1(new_n754), .B2(G128), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n765), .A2(G50), .B1(new_n753), .B2(G137), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1159), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n792), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n750), .B1(new_n274), .B2(new_n848), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1153), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1151), .A2(new_n1152), .A3(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n293), .A2(new_n869), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n305), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n305), .A2(new_n1175), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OR3_X1    g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n744), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n848), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n740), .B1(new_n1185), .B2(G50), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n753), .A2(G97), .B1(new_n827), .B2(new_n342), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT120), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n765), .A2(G58), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT119), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n309), .A2(G41), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n787), .B2(new_n757), .C1(new_n553), .C2(new_n773), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1054), .B1(new_n379), .B2(new_n767), .C1(new_n441), .C2(new_n829), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1188), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1191), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n280), .C1(G33), .C2(G41), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n773), .A2(new_n1199), .B1(new_n771), .B2(new_n830), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G132), .B2(new_n753), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G150), .A2(new_n768), .B1(new_n754), .B2(G125), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1163), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1202), .C1(new_n1203), .C2(new_n762), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n765), .A2(G159), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1198), .B1(KEYINPUT58), .B2(new_n1194), .C1(new_n1205), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1186), .B1(new_n1210), .B2(new_n792), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1184), .A2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT121), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n905), .A2(new_n928), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n678), .B1(new_n934), .B2(new_n906), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1182), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT122), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1218), .B1(new_n950), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1214), .A2(new_n1215), .A3(new_n1183), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1217), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1214), .A2(new_n1215), .A3(new_n1183), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1183), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT123), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1226), .B2(new_n950), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1213), .B1(new_n1227), .B2(new_n739), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1134), .A2(new_n1138), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1147), .B1(new_n1130), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1223), .A2(new_n1224), .B1(KEYINPUT124), .B2(new_n951), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n950), .B(KEYINPUT124), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1230), .A3(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n691), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1228), .B1(new_n1231), .B2(new_n1237), .ZN(G375));
  INV_X1    g1038(.A(new_n995), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1229), .A2(new_n1146), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1149), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n947), .A2(new_n744), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n740), .B1(new_n1185), .B2(G68), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n441), .A2(new_n831), .B1(new_n829), .B2(new_n788), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G97), .B2(new_n1021), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n771), .A2(new_n553), .B1(new_n757), .B2(new_n785), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n309), .B(new_n1246), .C1(G283), .C2(new_n776), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n1015), .A3(new_n1055), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n829), .A2(new_n837), .B1(new_n1057), .B2(new_n762), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G50), .B2(new_n768), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n771), .A2(new_n276), .B1(new_n757), .B2(new_n1199), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n259), .B(new_n1251), .C1(G137), .C2(new_n776), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(new_n831), .C2(new_n1203), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1248), .B1(new_n1253), .B2(new_n1190), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1243), .B1(new_n1254), .B2(new_n792), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1144), .A2(new_n739), .B1(new_n1242), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1241), .A2(new_n1256), .ZN(G381));
  OAI21_X1  g1057(.A(new_n1105), .B1(new_n1076), .B2(new_n738), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(G381), .ZN(new_n1263));
  OR4_X1    g1063(.A1(G387), .A2(new_n1263), .A3(G375), .A4(G378), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n1152), .A2(new_n1173), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n669), .A2(G213), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT125), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  OAI211_X1 g1070(.A(G378), .B(new_n1228), .C1(new_n1231), .C2(new_n1237), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1235), .A2(new_n739), .B1(new_n1184), .B2(new_n1211), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1222), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1219), .B1(new_n1233), .B2(new_n1218), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1230), .C1(new_n1274), .C2(new_n951), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1272), .B1(new_n1275), .B2(new_n995), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1266), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1271), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1139), .A2(new_n1143), .A3(KEYINPUT60), .A4(new_n1146), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n691), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT60), .B1(new_n1229), .B2(new_n1146), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1240), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1256), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1260), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1281), .A2(new_n1240), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G384), .B(new_n1256), .C1(new_n1285), .C2(new_n1280), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1278), .A2(new_n1267), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1278), .A2(new_n1267), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n669), .A2(G213), .A3(G2897), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1284), .A2(new_n1286), .A3(new_n1292), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1284), .A2(new_n1286), .B1(G2897), .B2(new_n1268), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(new_n809), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G390), .B(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1011), .A2(new_n1300), .A3(new_n1035), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1300), .B1(new_n1011), .B2(new_n1035), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1298), .B(new_n1259), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1011), .A2(new_n1300), .A3(new_n1035), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1303), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1268), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1290), .A2(new_n1297), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1308), .B1(new_n1310), .B2(new_n1295), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1288), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1310), .A2(KEYINPUT62), .A3(new_n1287), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1312), .B1(new_n1317), .B2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1266), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1271), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(KEYINPUT127), .A3(new_n1287), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1321), .A2(new_n1324), .A3(new_n1271), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1318), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1323), .A2(new_n1319), .A3(new_n1325), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


