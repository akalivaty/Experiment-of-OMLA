//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G567), .B1(G2106), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G113), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G113), .A3(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n467), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n472), .B2(G2105), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n459), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(G2105), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n475), .B1(new_n480), .B2(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(KEYINPUT4), .A2(G138), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n477), .B2(new_n478), .ZN(new_n487));
  AND2_X1   g062(.A1(G102), .A2(G2104), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n459), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  AND2_X1   g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G651), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n503), .B1(new_n500), .B2(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(G50), .A3(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(new_n510), .B1(new_n507), .B2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(new_n504), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n502), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(G63), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n511), .A2(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n504), .A3(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n504), .A2(G51), .A3(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT70), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n504), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n512), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n502), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n507), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n510), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT69), .B1(new_n509), .B2(KEYINPUT5), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n502), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(new_n546), .B2(new_n545), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n511), .A2(new_n504), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n504), .A2(G543), .ZN(new_n550));
  AOI22_X1  g125(.A1(G81), .A2(new_n549), .B1(new_n550), .B2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT72), .Z(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n543), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n549), .B2(G91), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n532), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n504), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND2_X1  g146(.A1(new_n549), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n550), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  OAI211_X1 g150(.A(G61), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n549), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n501), .A2(new_n503), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n500), .A2(G651), .ZN(new_n582));
  AND2_X1   g157(.A1(G48), .A2(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n504), .A2(KEYINPUT73), .A3(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n579), .A2(new_n580), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n543), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n502), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(new_n592), .ZN(new_n595));
  AOI22_X1  g170(.A1(G85), .A2(new_n549), .B1(new_n550), .B2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT75), .B1(new_n512), .B2(new_n599), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n543), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(new_n550), .B2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(G286), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(G299), .B(KEYINPUT76), .Z(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G297));
  AOI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g198(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  XOR2_X1   g201(.A(KEYINPUT77), .B(G2100), .Z(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n630), .B1(new_n480), .B2(new_n631), .C1(new_n632), .C2(new_n483), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n626), .A2(new_n627), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n628), .A2(new_n634), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(new_n653), .ZN(new_n660));
  INV_X1    g235(.A(new_n654), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n656), .A3(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(new_n655), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n658), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT79), .ZN(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n669), .A2(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n673), .A3(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n673), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT80), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  INV_X1    g260(.A(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n684), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n684), .B2(new_n688), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G23), .B(G288), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G1971), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n695), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT83), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  MUX2_X1   g282(.A(G24), .B(G290), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT81), .Z(new_n712));
  INV_X1    g287(.A(new_n483), .ZN(new_n713));
  INV_X1    g288(.A(new_n480), .ZN(new_n714));
  AOI22_X1  g289(.A1(G119), .A2(new_n713), .B1(new_n714), .B2(G131), .ZN(new_n715));
  NOR2_X1   g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT82), .Z(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n712), .B1(new_n719), .B2(G29), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n709), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n706), .A2(new_n707), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT36), .ZN(new_n725));
  AND3_X1   g300(.A1(G168), .A2(KEYINPUT90), .A3(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(KEYINPUT90), .B1(G168), .B2(G16), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G16), .B2(G21), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1966), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n699), .A2(G19), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n553), .B2(new_n699), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1341), .Z(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(KEYINPUT24), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(KEYINPUT24), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(KEYINPUT87), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT87), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G160), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n710), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n699), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n699), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n713), .A2(G129), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT88), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT26), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n746), .B(new_n748), .C1(new_n714), .C2(G141), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n710), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n710), .B2(G32), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT89), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n741), .B1(G1961), .B2(new_n743), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n710), .A2(G35), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n710), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G2090), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G11), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT30), .B(G28), .Z(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G29), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n633), .A2(new_n710), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(KEYINPUT91), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(KEYINPUT91), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n739), .A2(new_n740), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n710), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  INV_X1    g348(.A(G128), .ZN(new_n774));
  INV_X1    g349(.A(G140), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n774), .A2(new_n483), .B1(new_n480), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT84), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n466), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n776), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n773), .B1(new_n781), .B2(new_n710), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n752), .B2(new_n754), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n763), .A2(new_n771), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n756), .A2(new_n762), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n699), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n610), .B2(new_n699), .ZN(new_n788));
  INV_X1    g363(.A(G1348), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT95), .B(KEYINPUT23), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n699), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G299), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n699), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT96), .B(G1956), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n714), .A2(G139), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT86), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT85), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT25), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n802), .C1(new_n459), .C2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G33), .B(new_n804), .S(G29), .Z(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G2072), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n743), .A2(G1961), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT92), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n710), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n710), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2078), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n759), .B2(G2090), .ZN(new_n812));
  AND4_X1   g387(.A1(new_n797), .A2(new_n806), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n732), .A2(new_n786), .A3(new_n790), .A4(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n725), .A2(new_n729), .A3(new_n814), .ZN(G311));
  NAND3_X1  g390(.A1(new_n725), .A2(new_n729), .A3(new_n814), .ZN(G150));
  NAND2_X1  g391(.A1(new_n610), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  AOI22_X1  g393(.A1(G93), .A2(new_n549), .B1(new_n550), .B2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n502), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n552), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n818), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(G860), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n821), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(KEYINPUT100), .B(G37), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n781), .B(new_n497), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(new_n750), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n804), .A2(KEYINPUT98), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n750), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n804), .A2(KEYINPUT98), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n719), .B(KEYINPUT99), .ZN(new_n839));
  INV_X1    g414(.A(new_n625), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n714), .A2(G142), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n713), .A2(G130), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n839), .A2(new_n840), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n842), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n842), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n838), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n838), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(G160), .B(KEYINPUT97), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n633), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n853), .A2(new_n860), .A3(new_n854), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n831), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g438(.A(new_n620), .B(new_n822), .ZN(new_n864));
  INV_X1    g439(.A(new_n603), .ZN(new_n865));
  INV_X1    g440(.A(new_n609), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G299), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n610), .A2(new_n794), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(KEYINPUT41), .A3(new_n869), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n864), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G290), .B(G305), .ZN(new_n882));
  XNOR2_X1  g457(.A(G288), .B(G166), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n878), .A2(new_n886), .A3(new_n880), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(G868), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n885), .A2(new_n890), .A3(G868), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n821), .A2(new_n613), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(G295));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(G331));
  XOR2_X1   g469(.A(G168), .B(G301), .Z(new_n895));
  AND2_X1   g470(.A1(new_n822), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n822), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n871), .B2(new_n872), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n822), .B(new_n895), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n868), .B2(new_n869), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n884), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n872), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n903), .B2(new_n870), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n876), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n886), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n831), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n906), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n886), .B1(new_n904), .B2(new_n905), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n830), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT103), .B1(new_n913), .B2(KEYINPUT43), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n909), .B(new_n916), .C1(new_n911), .C2(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT102), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n902), .A2(new_n906), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n909), .A4(new_n916), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(KEYINPUT44), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n909), .B1(new_n919), .B2(new_n916), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI22_X1  g500(.A1(new_n915), .A2(new_n922), .B1(new_n925), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g501(.A1(new_n472), .A2(G2105), .ZN(new_n927));
  INV_X1    g502(.A(new_n464), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(G40), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n497), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT104), .Z(new_n935));
  INV_X1    g510(.A(new_n721), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n719), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n781), .B(G2067), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n750), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n934), .A2(G1996), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n750), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n938), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(G290), .A2(G1986), .A3(new_n934), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n949));
  AOI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n943), .B(KEYINPUT46), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n939), .A2(new_n750), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n935), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  INV_X1    g531(.A(G2067), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n781), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n942), .A2(new_n944), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n719), .A2(new_n936), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n935), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n951), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT124), .ZN(new_n964));
  INV_X1    g539(.A(new_n934), .ZN(new_n965));
  XNOR2_X1  g540(.A(G290), .B(G1986), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n945), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n929), .B1(new_n933), .B2(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(G2090), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n497), .A2(new_n971), .A3(new_n932), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT105), .B(G1971), .Z(new_n974));
  AOI21_X1  g549(.A(new_n929), .B1(new_n933), .B2(new_n931), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(G8), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G8), .B1(new_n514), .B2(new_n517), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT55), .B(G8), .C1(new_n514), .C2(new_n517), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n968), .B1(new_n978), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n933), .A2(new_n931), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(new_n930), .A3(new_n976), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n933), .A2(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(new_n930), .A3(new_n972), .ZN(new_n993));
  OAI22_X1  g568(.A1(new_n991), .A2(new_n974), .B1(G2090), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n984), .A2(new_n986), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n982), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT107), .A4(G8), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n988), .A2(new_n997), .B1(new_n978), .B2(new_n987), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n933), .A2(new_n929), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(G288), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT52), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1001), .B(new_n1005), .C1(new_n1002), .C2(G288), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  AOI22_X1  g586(.A1(G86), .A2(new_n549), .B1(new_n586), .B2(new_n587), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(new_n579), .ZN(new_n1013));
  AND4_X1   g588(.A1(new_n1011), .A2(new_n579), .A3(new_n580), .A4(new_n588), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1009), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1001), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1011), .A3(new_n579), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1010), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1008), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT49), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(KEYINPUT109), .A3(new_n1001), .A4(new_n1015), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1007), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n998), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n990), .B2(G2078), .ZN(new_n1028));
  INV_X1    g603(.A(G2078), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n975), .A2(KEYINPUT53), .A3(new_n1029), .A4(new_n976), .ZN(new_n1030));
  INV_X1    g605(.A(G1961), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n993), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1028), .A2(G301), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT122), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT123), .B1(new_n1035), .B2(G171), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1034), .B(KEYINPUT54), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1035), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT121), .B1(new_n1035), .B2(G171), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1033), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n993), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1044), .A2(new_n740), .B1(new_n990), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n528), .A2(G8), .A3(new_n529), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT119), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n990), .A2(new_n1045), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n969), .A2(new_n740), .A3(new_n972), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1000), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1047), .B(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1051), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n1058));
  OAI211_X1 g633(.A(new_n1048), .B(new_n1058), .C1(new_n1046), .C2(new_n1000), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1050), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1026), .A2(new_n1038), .A3(new_n1043), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1956), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n993), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n563), .A2(new_n568), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n975), .A2(new_n976), .A3(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1070));
  AND4_X1   g645(.A1(new_n930), .A2(new_n989), .A3(new_n976), .A4(new_n1067), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1956), .B1(new_n969), .B2(new_n972), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(KEYINPUT61), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1069), .B(new_n1073), .C1(KEYINPUT116), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n497), .A2(G160), .A3(G40), .A4(new_n932), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  AND3_X1   g656(.A1(new_n1080), .A2(KEYINPUT113), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT113), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n989), .A2(new_n940), .A3(new_n930), .A4(new_n976), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n975), .A2(KEYINPUT112), .A3(new_n940), .A4(new_n976), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n552), .B1(new_n1090), .B2(KEYINPUT59), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1090), .A2(KEYINPUT59), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n1093), .B(KEYINPUT115), .Z(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1089), .A2(new_n1094), .A3(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1079), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1079), .A2(KEYINPUT117), .A3(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n610), .A2(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n603), .B2(new_n609), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n993), .A2(new_n789), .B1(new_n957), .B2(new_n999), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT60), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n867), .A3(new_n1104), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1101), .A2(new_n1102), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n867), .A2(new_n1106), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1073), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1069), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1061), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n988), .A2(new_n997), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n978), .A2(new_n987), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1054), .A2(G168), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1025), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n998), .A2(new_n1025), .A3(KEYINPUT63), .A4(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1050), .A2(new_n1057), .A3(new_n1059), .A4(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1026), .A2(new_n1125), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1001), .B(KEYINPUT110), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G288), .A2(G1976), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1133), .B2(new_n1014), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT111), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1025), .A2(new_n988), .A3(new_n997), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1124), .B(new_n1129), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n964), .B(new_n967), .C1(new_n1116), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT111), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1125), .A2(new_n998), .A3(new_n1025), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1115), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1111), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1151), .B2(new_n1102), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1145), .B(new_n1148), .C1(new_n1152), .C2(new_n1061), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n964), .B1(new_n1153), .B2(new_n967), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n963), .B1(new_n1141), .B2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(G319), .ZN(new_n1157));
  NOR3_X1   g731(.A1(G401), .A2(new_n1157), .A3(G227), .ZN(new_n1158));
  OAI21_X1  g732(.A(new_n1158), .B1(new_n690), .B2(new_n691), .ZN(new_n1159));
  NOR3_X1   g733(.A1(new_n925), .A2(new_n862), .A3(new_n1159), .ZN(G308));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n862), .ZN(new_n1161));
  OAI21_X1  g735(.A(new_n1161), .B1(new_n924), .B2(new_n923), .ZN(G225));
endmodule


