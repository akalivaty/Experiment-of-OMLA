//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G15gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT28), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT27), .B1(new_n217), .B2(KEYINPUT66), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(G183gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT67), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n228), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n230), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n227), .A2(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT68), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n220), .A2(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n215), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT28), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT23), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n232), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT24), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT24), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n254), .A2(new_n256), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n217), .A2(new_n215), .ZN(new_n262));
  NAND3_X1  g061(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n253), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n225), .A2(new_n257), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n267), .A2(new_n262), .A3(new_n263), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n252), .B1(new_n268), .B2(new_n251), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G127gat), .A2(G134gat), .ZN(new_n271));
  INV_X1    g070(.A(G134gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G134gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n271), .B1(new_n276), .B2(G127gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G113gat), .B2(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G113gat), .ZN(new_n281));
  INV_X1    g080(.A(G120gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  NAND2_X1  g084(.A1(G127gat), .A2(G134gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n279), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n289));
  OAI21_X1  g088(.A(G113gat), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n246), .A2(new_n270), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n246), .B2(new_n270), .ZN(new_n294));
  NAND2_X1  g093(.A1(G227gat), .A2(G233gat), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n212), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n293), .B2(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT34), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT34), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n295), .C1(new_n293), .C2(new_n294), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n246), .A2(new_n270), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n277), .A2(new_n283), .B1(new_n287), .B2(new_n290), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n295), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n246), .A2(new_n270), .A3(new_n292), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n211), .B1(new_n310), .B2(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n309), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n302), .B1(new_n312), .B2(new_n295), .ZN(new_n313));
  INV_X1    g112(.A(new_n303), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(KEYINPUT32), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n304), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G78gat), .B(G106gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(G22gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT31), .B(G50gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G162gat), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G155gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  AND2_X1   g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT74), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(new_n341), .A3(new_n329), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n333), .A2(G155gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n331), .A2(G162gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT75), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n337), .A2(new_n340), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT76), .B(G155gat), .Z(new_n347));
  AOI21_X1  g146(.A(new_n328), .B1(new_n347), .B2(G162gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n335), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352));
  OR2_X1    g151(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n353));
  NAND2_X1  g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n356), .B2(new_n358), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT77), .B(new_n335), .C1(new_n346), .C2(new_n348), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n351), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n362), .B(new_n335), .C1(new_n346), .C2(new_n348), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n352), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n359), .A2(new_n360), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n368), .B1(new_n366), .B2(new_n352), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n340), .A2(new_n342), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT76), .B(G155gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT2), .B1(new_n377), .B2(new_n333), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n376), .A2(new_n378), .A3(new_n337), .A4(new_n345), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n362), .A2(new_n361), .B1(new_n379), .B2(new_n335), .ZN(new_n380));
  OR3_X1    g179(.A1(new_n375), .A2(new_n380), .A3(new_n373), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n324), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n365), .B2(new_n370), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n375), .A2(new_n380), .A3(new_n373), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n383), .A2(new_n384), .A3(new_n323), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n322), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n374), .A2(new_n381), .A3(new_n324), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n323), .B1(new_n383), .B2(new_n384), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n321), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n317), .B1(new_n304), .B2(new_n315), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n319), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n351), .A2(KEYINPUT3), .A3(new_n364), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n366), .A2(new_n292), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT4), .B1(new_n349), .B2(new_n292), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n379), .A2(new_n306), .A3(new_n398), .A4(new_n335), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n395), .A2(KEYINPUT5), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n396), .ZN(new_n402));
  AOI221_X4 g201(.A(new_n402), .B1(new_n397), .B2(new_n399), .C1(new_n393), .C2(new_n394), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n351), .A2(new_n364), .A3(new_n292), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n379), .A2(new_n335), .A3(new_n306), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n407), .B2(new_n402), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n401), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT0), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT6), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n396), .B1(new_n405), .B2(new_n406), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n416), .A2(new_n402), .B1(new_n417), .B2(new_n404), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n413), .A4(new_n401), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n413), .B(new_n401), .C1(new_n403), .C2(new_n408), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n243), .B1(new_n242), .B2(new_n244), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n433));
  OAI22_X1  g232(.A1(new_n236), .A2(KEYINPUT68), .B1(new_n433), .B2(new_n247), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n231), .A2(new_n227), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n225), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n437), .A2(new_n245), .B1(new_n269), .B2(new_n266), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n431), .B1(new_n246), .B2(new_n270), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n368), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n431), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n305), .B2(new_n352), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n444), .A2(new_n369), .A3(new_n440), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n430), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n369), .B1(new_n444), .B2(new_n440), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n246), .B2(new_n270), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n441), .B(new_n368), .C1(new_n443), .C2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n449), .A3(new_n429), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(KEYINPUT30), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n447), .A2(new_n449), .A3(new_n452), .A4(new_n429), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n392), .A2(new_n426), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n407), .A2(new_n402), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n393), .A2(new_n394), .B1(new_n397), .B2(new_n399), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n457), .A2(KEYINPUT5), .B1(new_n458), .B2(new_n396), .ZN(new_n459));
  INV_X1    g258(.A(new_n401), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n414), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n424), .A3(new_n421), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n425), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n386), .A2(new_n389), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n304), .A2(new_n315), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n316), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n466), .A2(new_n468), .A3(new_n454), .A4(new_n318), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n456), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n405), .A2(new_n406), .A3(new_n396), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT39), .B(new_n472), .C1(new_n458), .C2(new_n396), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n416), .A2(new_n474), .A3(new_n402), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT40), .A4(new_n414), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n421), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n396), .B1(new_n395), .B2(new_n400), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n413), .B1(new_n478), .B2(new_n474), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT40), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n454), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n390), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n442), .B2(new_n445), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n447), .A2(new_n449), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n430), .A4(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n488), .A2(new_n450), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n430), .A3(new_n487), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT38), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n489), .A2(new_n425), .A3(new_n462), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n468), .A2(KEYINPUT36), .A3(new_n318), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n319), .B2(new_n391), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n483), .A2(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n426), .A2(new_n454), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n390), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT79), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT79), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n471), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(G1gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(KEYINPUT83), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n505), .A2(G1gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(KEYINPUT83), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT84), .B(G8gat), .Z(new_n511));
  NAND4_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G8gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n209), .A2(G50gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n209), .A2(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT15), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n520), .B(KEYINPUT82), .Z(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n519), .A3(new_n525), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT80), .B(KEYINPUT15), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT81), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n522), .B1(new_n529), .B2(new_n524), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n209), .A2(KEYINPUT81), .A3(G50gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n521), .A2(new_n525), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n533), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT86), .B1(new_n515), .B2(new_n533), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(new_n538), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(new_n537), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n539), .A2(new_n540), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT11), .B(G169gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n541), .A2(new_n546), .A3(new_n553), .A4(new_n547), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT87), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n504), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n426), .ZN(new_n561));
  XOR2_X1   g360(.A(G57gat), .B(G64gat), .Z(new_n562));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g363(.A(G71gat), .ZN(new_n565));
  INV_X1    g364(.A(G78gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n562), .A2(new_n563), .A3(new_n569), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G127gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n516), .B1(new_n574), .B2(new_n573), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT89), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n331), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n586), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G99gat), .ZN(new_n590));
  INV_X1    g389(.A(G106gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT91), .B(KEYINPUT7), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(G85gat), .A3(G92gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n592), .A2(new_n594), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(new_n593), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n600), .B(new_n602), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n606), .A2(new_n593), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n599), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n608), .B(new_n611), .C1(new_n534), .C2(new_n535), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n611), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n613), .A2(new_n533), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT90), .ZN(new_n622));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n618), .B2(new_n619), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n573), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n605), .A2(new_n607), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n610), .B1(new_n609), .B2(new_n599), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n608), .A2(new_n611), .A3(new_n573), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n632), .B1(new_n641), .B2(KEYINPUT93), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n643), .A3(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n636), .A2(new_n638), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n632), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n641), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n631), .B(KEYINPUT94), .Z(new_n653));
  OAI21_X1  g452(.A(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n630), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n560), .A2(new_n561), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n560), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(G8gat), .B1(new_n661), .B2(new_n454), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT96), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n454), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  AOI21_X1  g464(.A(KEYINPUT95), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(G1325gat));
  NOR2_X1   g468(.A1(new_n319), .A2(new_n391), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n207), .B1(new_n661), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT97), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n495), .A2(new_n493), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n661), .A2(new_n207), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n466), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n589), .ZN(new_n680));
  INV_X1    g479(.A(new_n657), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n629), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n504), .A2(new_n559), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n426), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT45), .Z(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n629), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n501), .A2(new_n503), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n557), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT99), .B1(new_n456), .B2(new_n470), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n423), .A2(new_n425), .B1(new_n453), .B2(new_n451), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n464), .B1(new_n693), .B2(new_n392), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n465), .A2(new_n469), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n491), .A2(new_n450), .A3(new_n488), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n463), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n473), .A2(new_n475), .A3(new_n414), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n421), .A3(new_n476), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n466), .B1(new_n704), .B2(new_n454), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n674), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n693), .A2(new_n466), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT98), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT98), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n496), .A2(new_n709), .A3(new_n498), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n629), .B1(new_n698), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n689), .B(new_n691), .C1(new_n712), .C2(KEYINPUT44), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n706), .A2(KEYINPUT98), .A3(new_n707), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n709), .B1(new_n496), .B2(new_n498), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n456), .A2(KEYINPUT99), .A3(new_n470), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n696), .B1(new_n694), .B2(new_n695), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n628), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n687), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n723), .A2(KEYINPUT100), .A3(new_n689), .A4(new_n691), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n715), .A2(new_n724), .A3(new_n561), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G29gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n686), .A2(new_n726), .ZN(G1328gat));
  OR2_X1    g526(.A1(new_n454), .A2(G36gat), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n684), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n724), .A3(new_n482), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G36gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1329gat));
  NAND4_X1  g534(.A1(new_n560), .A2(new_n209), .A3(new_n670), .A4(new_n683), .ZN(new_n736));
  OAI21_X1  g535(.A(G43gat), .B1(new_n713), .B2(new_n674), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT47), .ZN(new_n738));
  INV_X1    g537(.A(new_n674), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n715), .A2(new_n724), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n736), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n738), .B1(new_n742), .B2(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g542(.A1(new_n466), .A2(G50gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n713), .B2(new_n466), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n713), .A2(new_n745), .A3(new_n466), .ZN(new_n748));
  OAI221_X1 g547(.A(KEYINPUT48), .B1(new_n684), .B2(new_n744), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n715), .A2(new_n724), .A3(new_n390), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n750), .A2(KEYINPUT102), .A3(G50gat), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT102), .B1(new_n750), .B2(G50gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n684), .A2(new_n744), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n749), .B1(new_n754), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g554(.A1(new_n718), .A2(new_n721), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n756), .A2(new_n557), .A3(new_n630), .A4(new_n681), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n561), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g558(.A(new_n454), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1333gat));
  AOI21_X1  g564(.A(new_n565), .B1(new_n757), .B2(new_n739), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n671), .A2(G71gat), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n757), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n390), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n589), .A2(new_n557), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT51), .B1(new_n712), .B2(new_n772), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n561), .A2(new_n596), .A3(new_n657), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n723), .A2(new_n657), .A3(new_n689), .A4(new_n772), .ZN(new_n781));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781), .B2(new_n426), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1336gat));
  NOR3_X1   g582(.A1(new_n681), .A2(G92gat), .A3(new_n454), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n781), .B2(new_n454), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n773), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n784), .B1(new_n789), .B2(new_n776), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n786), .B2(new_n791), .ZN(G1337gat));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n590), .A3(new_n670), .A4(new_n657), .ZN(new_n793));
  OAI21_X1  g592(.A(G99gat), .B1(new_n781), .B2(new_n674), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n657), .A2(new_n591), .A3(new_n390), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT108), .Z(new_n797));
  AOI21_X1  g596(.A(KEYINPUT53), .B1(new_n777), .B2(new_n797), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n466), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT111), .B1(new_n781), .B2(new_n466), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(G106gat), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n781), .B2(new_n466), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n797), .B(KEYINPUT109), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n789), .B2(new_n776), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n806), .B2(KEYINPUT53), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n806), .A2(KEYINPUT110), .A3(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n658), .A2(new_n690), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(KEYINPUT114), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n813), .B(new_n814), .C1(new_n545), .C2(new_n543), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n552), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n628), .A2(new_n816), .A3(new_n556), .ZN(new_n817));
  INV_X1    g616(.A(new_n653), .ZN(new_n818));
  XOR2_X1   g617(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n819));
  NAND3_X1  g618(.A1(new_n641), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n655), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n641), .A2(KEYINPUT93), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n823), .A2(new_n631), .A3(new_n644), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n639), .A2(new_n640), .A3(new_n653), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(KEYINPUT55), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n651), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n642), .B2(new_n644), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n821), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n830), .A3(new_n821), .ZN(new_n833));
  INV_X1    g632(.A(new_n651), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n817), .A2(new_n829), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n835), .A2(new_n557), .A3(new_n829), .A4(new_n832), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n816), .A2(new_n556), .A3(new_n657), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n628), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(KEYINPUT115), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n589), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n840), .A2(new_n841), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n629), .A3(new_n843), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n836), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT116), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n811), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n390), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(new_n561), .A3(new_n454), .A4(new_n670), .ZN(new_n853));
  OAI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n558), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n851), .A2(new_n426), .A3(new_n469), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n557), .A2(new_n281), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  OAI21_X1  g657(.A(G120gat), .B1(new_n853), .B2(new_n681), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n681), .A2(new_n288), .A3(new_n289), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n856), .B2(new_n860), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n853), .B2(new_n680), .ZN(new_n862));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n855), .A2(new_n863), .A3(new_n589), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1342gat));
  NOR2_X1   g664(.A1(new_n851), .A2(new_n426), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n629), .A2(new_n276), .A3(new_n482), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n392), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT56), .Z(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n853), .B2(new_n629), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  NAND3_X1  g670(.A1(new_n848), .A2(new_n845), .A3(new_n836), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n680), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n844), .A2(new_n845), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n810), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n390), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n739), .A2(new_n426), .A3(new_n482), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n827), .A2(new_n832), .A3(new_n651), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n558), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n839), .B(KEYINPUT118), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n629), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n589), .B1(new_n883), .B2(new_n836), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n390), .B1(new_n884), .B2(new_n811), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n879), .B1(new_n885), .B2(KEYINPUT57), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n325), .B1(new_n887), .B2(new_n557), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n739), .A2(new_n466), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n482), .ZN(new_n891));
  AND4_X1   g690(.A1(new_n325), .A2(new_n866), .A3(new_n559), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n559), .A3(new_n886), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n877), .A2(new_n886), .A3(KEYINPUT119), .A4(new_n559), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(G141gat), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n900), .ZN(G1344gat));
  NAND4_X1  g700(.A1(new_n866), .A2(new_n326), .A3(new_n657), .A4(new_n891), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n875), .A2(new_n390), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n559), .A2(new_n630), .A3(new_n657), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n884), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n466), .A2(KEYINPUT57), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n906), .A2(KEYINPUT57), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n657), .A3(new_n878), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n905), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT59), .B(new_n326), .C1(new_n887), .C2(new_n657), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(G1345gat));
  AND2_X1   g713(.A1(new_n866), .A2(new_n891), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n377), .A3(new_n589), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n877), .A2(new_n886), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n347), .B1(new_n917), .B2(new_n680), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1346gat));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n333), .A3(new_n628), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n917), .B2(new_n629), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G162gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n917), .A2(new_n921), .A3(new_n629), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n851), .A2(new_n561), .ZN(new_n926));
  INV_X1    g725(.A(new_n392), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n454), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n557), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n561), .A2(new_n454), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n671), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n852), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n229), .A3(new_n558), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n930), .A2(new_n935), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n230), .A3(new_n657), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n934), .B2(new_n681), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  NAND4_X1  g738(.A1(new_n926), .A2(new_n214), .A3(new_n589), .A4(new_n928), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n934), .A2(new_n680), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n217), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI221_X1 g744(.A(new_n940), .B1(KEYINPUT122), .B2(new_n943), .C1(new_n941), .C2(new_n217), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1350gat));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n629), .A2(G190gat), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n926), .A2(new_n948), .A3(new_n928), .A4(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n875), .A2(new_n426), .A3(new_n928), .A4(new_n949), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n875), .A2(new_n466), .A3(new_n628), .A4(new_n933), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G190gat), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n953), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n953), .A2(new_n957), .A3(KEYINPUT124), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1351gat));
  NOR4_X1   g762(.A1(new_n851), .A2(new_n561), .A3(new_n454), .A4(new_n890), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n557), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n932), .A2(new_n739), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n910), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n559), .A2(G197gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  NAND3_X1  g768(.A1(new_n910), .A2(new_n657), .A3(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G204gat), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n681), .A2(G204gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT62), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n971), .B(new_n974), .C1(new_n976), .C2(new_n977), .ZN(G1353gat));
  INV_X1    g777(.A(G211gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n979), .A3(new_n589), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT57), .B1(new_n851), .B2(new_n466), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n908), .A2(new_n909), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n981), .A2(new_n589), .A3(new_n982), .A4(new_n966), .ZN(new_n983));
  AND4_X1   g782(.A1(KEYINPUT126), .A2(new_n983), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AOI22_X1  g785(.A1(new_n983), .A2(new_n986), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n980), .B1(new_n984), .B2(new_n987), .ZN(G1354gat));
  AOI21_X1  g787(.A(KEYINPUT127), .B1(new_n910), .B2(new_n966), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n981), .A2(KEYINPUT127), .A3(new_n982), .A4(new_n966), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n628), .ZN(new_n991));
  OAI21_X1  g790(.A(G218gat), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(G218gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n964), .A2(new_n993), .A3(new_n628), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1355gat));
endmodule


