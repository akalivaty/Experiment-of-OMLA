//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G227), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G146), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n193), .A2(KEYINPUT65), .A3(G143), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n194), .B(new_n196), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT82), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n194), .B1(new_n199), .B2(new_n200), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g019(.A(G128), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(KEYINPUT83), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT65), .B1(new_n193), .B2(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n197), .A2(new_n198), .A3(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n195), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n214), .A3(new_n196), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n202), .A2(new_n207), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G104), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n222), .A2(new_n228), .A3(G101), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT81), .ZN(new_n230));
  XNOR2_X1  g044(.A(G104), .B(G107), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n223), .A2(G104), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT81), .B(G101), .C1(new_n219), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT10), .B1(new_n216), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n198), .A3(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n194), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n244), .A2(new_n246), .B1(new_n211), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(G101), .C1(new_n222), .C2(new_n228), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(G101), .B1(new_n222), .B2(new_n228), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n234), .B1(new_n224), .B2(new_n226), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n219), .B1(new_n221), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n256), .A3(new_n232), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n257), .A3(KEYINPUT4), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n244), .A2(new_n206), .B1(new_n211), .B2(new_n196), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT10), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n252), .A2(new_n258), .B1(new_n261), .B2(new_n237), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT66), .A2(G137), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT66), .A2(G137), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT11), .A2(G134), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G131), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT11), .A2(G134), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT11), .A2(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(new_n266), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n239), .A2(new_n262), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n216), .A2(new_n237), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n257), .A2(new_n235), .A3(new_n233), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n259), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n270), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n270), .A3(new_n267), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT12), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n284), .B(new_n273), .C1(new_n275), .C2(new_n277), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n192), .B(new_n274), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n273), .B1(new_n239), .B2(new_n262), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n253), .A2(new_n257), .A3(KEYINPUT4), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n249), .A2(new_n251), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n204), .B1(new_n240), .B2(new_n242), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n201), .B1(new_n290), .B2(new_n212), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n288), .A2(new_n289), .B1(new_n292), .B2(new_n276), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n293), .A2(new_n238), .A3(new_n282), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n191), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT71), .B(G902), .Z(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n294), .A2(new_n191), .ZN(new_n300));
  INV_X1    g114(.A(new_n287), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n278), .A2(new_n282), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n284), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n278), .A2(KEYINPUT12), .A3(new_n282), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n302), .B(G469), .C1(new_n306), .C2(new_n192), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n297), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n299), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G221), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n298), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n286), .B2(new_n295), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n309), .B1(new_n321), .B2(new_n297), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n322), .B2(new_n307), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT84), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n232), .B1(new_n254), .B2(new_n256), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n329));
  INV_X1    g143(.A(G113), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT2), .A2(G113), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G116), .B(G119), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n331), .A2(new_n332), .B1(KEYINPUT2), .B2(G113), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n336), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n327), .A2(new_n250), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G116), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G119), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n330), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G116), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(G119), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT5), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n339), .A2(new_n336), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n341), .A2(new_n258), .B1(new_n237), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G122), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n326), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n352), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n351), .B2(KEYINPUT85), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n350), .A2(new_n257), .A3(new_n235), .A4(new_n233), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n339), .A2(new_n336), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n251), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n288), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n244), .A2(new_n206), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(new_n201), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n247), .B(new_n204), .C1(new_n209), .C2(new_n210), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n245), .B1(new_n243), .B2(new_n194), .ZN(new_n369));
  OAI21_X1  g183(.A(G125), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n365), .B1(new_n259), .B2(new_n366), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G953), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G224), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT87), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n373), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n351), .A2(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n360), .A2(new_n361), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n326), .A4(new_n354), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n363), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n375), .A2(KEYINPUT7), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n382), .B(new_n383), .C1(new_n371), .C2(new_n372), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n356), .B(new_n352), .C1(new_n288), .C2(new_n359), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n350), .B1(new_n229), .B2(new_n236), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n352), .B(KEYINPUT8), .ZN(new_n388));
  OAI21_X1  g202(.A(G113), .B1(new_n347), .B2(KEYINPUT5), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n389), .A2(new_n390), .B1(new_n336), .B2(KEYINPUT5), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n345), .A2(KEYINPUT88), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n391), .A2(new_n392), .B1(new_n339), .B2(new_n336), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n387), .B(new_n388), .C1(new_n276), .C2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n201), .B(new_n366), .C1(new_n290), .C2(new_n212), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT86), .ZN(new_n396));
  INV_X1    g210(.A(new_n383), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n396), .A2(new_n370), .A3(new_n367), .A4(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n386), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n385), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT89), .B1(new_n373), .B2(new_n397), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G210), .B1(G237), .B2(G902), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n381), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n381), .A2(new_n402), .A3(KEYINPUT91), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n381), .A2(new_n402), .ZN(new_n409));
  INV_X1    g223(.A(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT90), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n403), .B1(new_n381), .B2(new_n402), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n408), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n217), .ZN(new_n418));
  INV_X1    g232(.A(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n366), .A2(G140), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(KEYINPUT75), .A3(G125), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT16), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G146), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n420), .A2(new_n421), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT19), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n193), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT69), .B(G237), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(G214), .A3(new_n374), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n198), .ZN(new_n437));
  OR2_X1    g251(.A1(KEYINPUT69), .A2(G237), .ZN(new_n438));
  NAND2_X1  g252(.A1(KEYINPUT69), .A2(G237), .ZN(new_n439));
  AOI21_X1  g253(.A(G953), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(G143), .A3(G214), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n267), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n267), .B1(new_n437), .B2(new_n441), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n429), .B(new_n434), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n437), .A2(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT18), .A3(G131), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n423), .A2(G146), .A3(new_n424), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n432), .A2(new_n193), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT18), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n437), .B(new_n441), .C1(new_n451), .C2(new_n267), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n418), .B1(new_n445), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n450), .ZN(new_n455));
  AOI211_X1 g269(.A(new_n451), .B(new_n267), .C1(new_n437), .C2(new_n441), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n425), .A2(new_n193), .A3(new_n427), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n429), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(KEYINPUT17), .B2(new_n444), .ZN(new_n460));
  INV_X1    g274(.A(new_n444), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT17), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n442), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n457), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n454), .B1(new_n464), .B2(new_n418), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT92), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT20), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n469));
  INV_X1    g283(.A(new_n467), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT17), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n446), .A2(KEYINPUT17), .A3(G131), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n429), .A3(new_n458), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n418), .B(new_n453), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n469), .B(new_n470), .C1(new_n475), .C2(new_n454), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n453), .B1(new_n471), .B2(new_n473), .ZN(new_n478));
  INV_X1    g292(.A(new_n418), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n480), .A2(new_n474), .ZN(new_n481));
  OAI21_X1  g295(.A(G475), .B1(new_n481), .B2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G122), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G116), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n342), .A2(G122), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n223), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT94), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n484), .A2(G116), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n485), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT95), .B1(new_n486), .B2(KEYINPUT14), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n497), .B(G107), .C1(new_n495), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G128), .B(G143), .ZN(new_n500));
  INV_X1    g314(.A(G134), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n342), .A2(G122), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT93), .B1(new_n503), .B2(new_n493), .ZN(new_n504));
  AOI21_X1  g318(.A(G107), .B1(new_n504), .B2(new_n488), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n492), .A2(new_n499), .A3(new_n502), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT13), .B1(new_n195), .B2(G143), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n501), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n500), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n489), .A2(new_n223), .A3(new_n490), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n505), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G217), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n313), .A2(new_n515), .A3(G953), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n513), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n298), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n320), .B1(new_n518), .B2(new_n519), .ZN(new_n526));
  INV_X1    g340(.A(new_n524), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT96), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n298), .A3(new_n527), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT97), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(KEYINPUT97), .A3(new_n527), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G952), .ZN(new_n536));
  AOI211_X1 g350(.A(G953), .B(new_n536), .C1(G234), .C2(G237), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n374), .B(new_n298), .C1(G234), .C2(G237), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT21), .B(G898), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT98), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n483), .A2(new_n535), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n416), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n187), .B1(new_n325), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n311), .A2(KEYINPUT84), .A3(new_n316), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT84), .B1(new_n311), .B2(new_n316), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n544), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n413), .A2(new_n414), .ZN(new_n551));
  AOI211_X1 g365(.A(KEYINPUT90), .B(new_n403), .C1(new_n381), .C2(new_n402), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n550), .B1(new_n553), .B2(new_n408), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n549), .A2(KEYINPUT99), .A3(new_n543), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n440), .A2(G210), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT27), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT27), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n440), .A2(new_n558), .A3(G210), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n263), .A2(new_n501), .A3(new_n264), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n267), .B1(G134), .B2(G137), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n281), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n291), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n244), .A2(new_n246), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n211), .A2(new_n248), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n573), .C1(new_n271), .C2(new_n272), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n357), .A2(new_n358), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n203), .A2(new_n247), .B1(new_n290), .B2(new_n245), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT67), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n273), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT67), .B1(new_n282), .B2(new_n249), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n571), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT30), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n571), .A2(new_n574), .A3(KEYINPUT30), .ZN(new_n585));
  INV_X1    g399(.A(new_n575), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n577), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n566), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n576), .A2(KEYINPUT28), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT28), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n249), .A2(new_n282), .B1(new_n570), .B2(new_n291), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n575), .ZN(new_n595));
  INV_X1    g409(.A(new_n571), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n574), .A2(new_n579), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n282), .A2(new_n249), .A3(KEYINPUT67), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n592), .A2(new_n595), .B1(new_n599), .B2(new_n575), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n563), .A2(KEYINPUT70), .A3(new_n564), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT70), .B1(new_n563), .B2(new_n564), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n590), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n594), .A2(new_n575), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n576), .A2(KEYINPUT28), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n594), .A2(new_n593), .A3(new_n575), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n600), .A2(new_n604), .B1(new_n608), .B2(new_n590), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n298), .B1(new_n591), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n587), .B1(new_n583), .B2(new_n582), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n566), .A2(new_n576), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT31), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT31), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n577), .A2(new_n565), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n599), .A2(KEYINPUT30), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n587), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n602), .A2(new_n603), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n614), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT32), .ZN(new_n622));
  NOR2_X1   g436(.A1(G472), .A2(G902), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n611), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT72), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT22), .B(G137), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n374), .A2(G221), .A3(G234), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n628), .B(new_n629), .Z(new_n630));
  OAI211_X1 g444(.A(new_n195), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT23), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n346), .B2(G128), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT73), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n346), .B2(G128), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G110), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT74), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT74), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n639), .A3(G110), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT24), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(G119), .B(G128), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n638), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT77), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT76), .B1(new_n641), .B2(new_n642), .ZN(new_n646));
  INV_X1    g460(.A(G110), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n647), .B(new_n631), .C1(new_n633), .C2(new_n635), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT24), .B(G110), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT76), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n346), .A2(G128), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n346), .A2(G128), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n649), .B(new_n650), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n646), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n449), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n193), .B1(new_n425), .B2(new_n427), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n645), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n429), .A2(KEYINPUT77), .A3(new_n655), .A4(new_n449), .ZN(new_n659));
  AOI221_X4 g473(.A(KEYINPUT78), .B1(new_n644), .B2(new_n459), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT78), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n644), .A2(new_n459), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n630), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n630), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(KEYINPUT78), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n298), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT25), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n665), .A2(KEYINPUT25), .A3(new_n298), .A4(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n515), .B1(new_n298), .B2(G234), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n665), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT79), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT79), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n665), .A2(new_n677), .A3(new_n668), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n674), .A2(G902), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n673), .A2(new_n674), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT72), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n611), .B(new_n682), .C1(new_n624), .C2(new_n625), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n627), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n546), .A2(new_n555), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT100), .B(G101), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G3));
  INV_X1    g501(.A(new_n681), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n621), .A2(new_n623), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n621), .A2(new_n298), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n689), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n549), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n477), .A2(new_n482), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n520), .B(KEYINPUT33), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n320), .A2(new_n523), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n699), .A2(new_n700), .B1(new_n523), .B2(new_n521), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n404), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n544), .B1(new_n703), .B2(new_n413), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n542), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n697), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT34), .B(G104), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G6));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n525), .A2(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n483), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n713), .B1(new_n716), .B2(new_n542), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(KEYINPUT104), .A3(new_n706), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n705), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n697), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT35), .B(G107), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G9));
  NOR2_X1   g536(.A1(new_n667), .A2(KEYINPUT105), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n662), .B2(new_n663), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n666), .A2(KEYINPUT36), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OR3_X1    g541(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n723), .B2(new_n725), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(new_n680), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n673), .B2(new_n674), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n695), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n546), .A2(new_n555), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT37), .B(G110), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G12));
  INV_X1    g549(.A(G900), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n537), .B1(new_n538), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n483), .A2(new_n714), .A3(new_n737), .ZN(new_n738));
  AND4_X1   g552(.A1(new_n319), .A2(new_n324), .A3(new_n705), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n673), .A2(new_n674), .ZN(new_n740));
  INV_X1    g554(.A(new_n730), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n627), .A2(new_n683), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G128), .ZN(G30));
  XOR2_X1   g559(.A(new_n737), .B(KEYINPUT39), .Z(new_n746));
  NAND2_X1  g560(.A1(new_n549), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT40), .Z(new_n748));
  XOR2_X1   g562(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n416), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(G472), .A2(G902), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n612), .A2(new_n613), .ZN(new_n752));
  INV_X1    g566(.A(new_n603), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n601), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n605), .A2(new_n577), .ZN(new_n755));
  OAI21_X1  g569(.A(G472), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n751), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT107), .Z(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n625), .B2(new_n624), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n483), .A2(new_n535), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n550), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n731), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n750), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n748), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G143), .ZN(G45));
  AND2_X1   g579(.A1(new_n627), .A2(new_n683), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n547), .A2(new_n731), .A3(new_n548), .ZN(new_n767));
  INV_X1    g581(.A(new_n701), .ZN(new_n768));
  INV_X1    g582(.A(new_n737), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n483), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n704), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G146), .ZN(G48));
  NAND3_X1  g587(.A1(new_n627), .A2(new_n681), .A3(new_n683), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n296), .A2(new_n298), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(G469), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n299), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT108), .A3(G469), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n316), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n774), .A2(new_n707), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT41), .B(G113), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G15));
  NOR3_X1   g598(.A1(new_n719), .A2(new_n774), .A3(new_n781), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n342), .ZN(G18));
  AOI21_X1  g600(.A(new_n315), .B1(new_n778), .B2(new_n779), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n543), .A3(new_n705), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n627), .A2(new_n742), .A3(new_n683), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n346), .ZN(G21));
  NOR3_X1   g605(.A1(new_n704), .A2(new_n760), .A3(new_n542), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n608), .A2(new_n754), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n614), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n614), .A3(KEYINPUT109), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n618), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n798), .A2(new_n623), .B1(G472), .B2(new_n690), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(new_n681), .A3(new_n787), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G122), .ZN(G24));
  NOR2_X1   g615(.A1(new_n781), .A2(new_n704), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n698), .A2(new_n701), .A3(new_n737), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n742), .A2(new_n803), .A3(new_n799), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT110), .B(G125), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G27));
  NAND4_X1  g621(.A1(new_n553), .A2(new_n323), .A3(new_n544), .A4(new_n408), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n681), .A2(new_n626), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT42), .A4(new_n803), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n684), .A2(KEYINPUT111), .A3(new_n803), .A4(new_n809), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT42), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n774), .A2(new_n808), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT111), .B1(new_n815), .B2(new_n803), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n811), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G131), .ZN(G33));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n738), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  NAND3_X1  g634(.A1(new_n553), .A2(new_n544), .A3(new_n408), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n698), .A2(new_n768), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT43), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n695), .A3(new_n742), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT44), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n302), .B1(new_n306), .B2(new_n192), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT45), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n297), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(KEYINPUT46), .A3(new_n310), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n829), .B1(new_n834), .B2(new_n299), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT46), .B1(new_n833), .B2(new_n310), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n829), .A3(new_n299), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n316), .A3(new_n746), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(G137), .Z(G39));
  AOI21_X1  g656(.A(new_n315), .B1(new_n837), .B2(new_n838), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT47), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(KEYINPUT47), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n766), .A2(new_n681), .A3(new_n770), .A4(new_n821), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G140), .ZN(G42));
  XNOR2_X1  g663(.A(new_n780), .B(KEYINPUT49), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n688), .A2(new_n759), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n822), .A2(new_n315), .A3(new_n550), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n750), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT113), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n702), .A2(new_n715), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n542), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n696), .A3(new_n549), .A4(new_n554), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n685), .A2(new_n733), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n800), .B1(new_n788), .B2(new_n789), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n785), .A2(new_n860), .A3(new_n782), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n815), .A2(new_n738), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n804), .A2(new_n809), .ZN(new_n863));
  INV_X1    g677(.A(new_n821), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n483), .A2(new_n535), .A3(new_n737), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n627), .A3(new_n683), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n767), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n817), .A2(new_n859), .A3(new_n861), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n317), .A2(new_n737), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n704), .A2(new_n760), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n759), .A2(new_n871), .A3(new_n872), .A4(new_n731), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n744), .A2(new_n772), .A3(new_n805), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n743), .A2(new_n739), .B1(new_n802), .B2(new_n804), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n772), .A4(new_n873), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n855), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n685), .A2(new_n733), .A3(new_n858), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n819), .B(new_n863), .C1(new_n867), .C2(new_n866), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n855), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n876), .A2(new_n878), .B1(KEYINPUT114), .B2(new_n874), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n874), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n811), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n774), .A2(new_n770), .A3(new_n808), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT42), .B1(new_n889), .B2(KEYINPUT111), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n684), .A2(new_n803), .A3(new_n809), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT111), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n860), .A2(new_n782), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n719), .A2(new_n774), .A3(new_n781), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT116), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n817), .A2(new_n899), .A3(new_n861), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n880), .B(new_n881), .C1(new_n887), .C2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT117), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n882), .A2(new_n883), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n876), .A2(new_n878), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n817), .A4(new_n861), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n855), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n874), .A2(KEYINPUT114), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n886), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n855), .B1(new_n909), .B2(new_n870), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(new_n910), .B2(KEYINPUT115), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n912), .B(new_n855), .C1(new_n909), .C2(new_n870), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n881), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n864), .A2(new_n537), .A3(new_n787), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n810), .A3(new_n824), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT48), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n536), .A2(G953), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n702), .A3(new_n851), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n824), .A2(new_n537), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n681), .A2(new_n799), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n802), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n915), .A2(new_n698), .A3(new_n701), .A4(new_n851), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n915), .A2(new_n742), .A3(new_n799), .A4(new_n824), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(KEYINPUT120), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n921), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT50), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n750), .A2(new_n550), .A3(new_n787), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n926), .A2(KEYINPUT120), .ZN(new_n934));
  AND4_X1   g748(.A1(KEYINPUT51), .A2(new_n927), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n780), .A2(new_n315), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n844), .A2(new_n845), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n920), .A2(new_n921), .A3(new_n864), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT118), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n923), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(KEYINPUT119), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT119), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n937), .B2(new_n939), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n933), .A2(new_n926), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n941), .B1(new_n946), .B2(KEYINPUT51), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n903), .A2(new_n914), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(G952), .A2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n854), .B1(new_n948), .B2(new_n949), .ZN(G75));
  OAI21_X1  g764(.A(new_n880), .B1(new_n887), .B2(new_n901), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n951), .A2(new_n320), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n410), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n363), .A2(new_n380), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT121), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n377), .B(KEYINPUT55), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n953), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n953), .B2(new_n954), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n374), .A2(G952), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G51));
  NAND2_X1  g776(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n964), .A3(new_n902), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n951), .A2(KEYINPUT122), .A3(KEYINPUT54), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n309), .B(KEYINPUT57), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n296), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n833), .B(KEYINPUT123), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n952), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n961), .B1(new_n969), .B2(new_n971), .ZN(G54));
  NAND3_X1  g786(.A1(new_n952), .A2(KEYINPUT58), .A3(G475), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(new_n465), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n465), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(new_n961), .ZN(G60));
  INV_X1    g790(.A(new_n699), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT59), .Z(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n965), .A2(new_n966), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n961), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n979), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n903), .B2(new_n914), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n977), .B2(new_n985), .ZN(G63));
  AND2_X1   g800(.A1(new_n728), .A2(new_n729), .ZN(new_n987));
  XNOR2_X1  g801(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n515), .A2(new_n308), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n951), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(KEYINPUT125), .A3(new_n982), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT61), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n951), .A2(new_n990), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n982), .B(new_n991), .C1(new_n994), .C2(new_n679), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G66));
  INV_X1    g810(.A(G224), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n541), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n897), .A2(new_n882), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n956), .B1(G898), .B2(new_n374), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  NAND2_X1  g816(.A1(new_n584), .A2(new_n585), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n431), .A2(new_n433), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n764), .A2(new_n772), .A3(new_n877), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  NOR4_X1   g822(.A1(new_n747), .A2(new_n774), .A3(new_n821), .A4(new_n856), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n841), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n764), .A2(new_n1011), .A3(new_n772), .A4(new_n877), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1008), .A2(new_n1010), .A3(new_n848), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1006), .B1(new_n1013), .B2(new_n374), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n894), .B1(new_n846), .B2(new_n847), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n843), .A2(new_n746), .A3(new_n872), .A4(new_n810), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n877), .A2(new_n772), .A3(new_n819), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n841), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n374), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(G900), .B2(new_n374), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1014), .B1(new_n1021), .B2(new_n1006), .ZN(new_n1022));
  OAI21_X1  g836(.A(G953), .B1(new_n189), .B2(new_n736), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT126), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1022), .B(new_n1024), .ZN(G72));
  XOR2_X1   g839(.A(new_n751), .B(KEYINPUT63), .Z(new_n1026));
  INV_X1    g840(.A(new_n999), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1026), .B1(new_n1013), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n589), .A2(new_n565), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n961), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1015), .A2(new_n999), .A3(new_n1018), .A4(new_n1016), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1031), .A2(new_n1032), .A3(new_n1026), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n612), .A2(new_n577), .A3(new_n566), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n1031), .B2(new_n1026), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1030), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n911), .A2(new_n913), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1026), .ZN(new_n1039));
  NOR3_X1   g853(.A1(new_n1029), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1037), .B1(new_n1038), .B2(new_n1040), .ZN(G57));
endmodule


