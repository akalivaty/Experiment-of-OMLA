//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n203));
  INV_X1    g002(.A(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT78), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G197gat), .ZN(new_n206));
  INV_X1    g005(.A(G197gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT78), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(KEYINPUT78), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(G197gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(G204gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n203), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g015(.A(KEYINPUT79), .B(new_n214), .C1(new_n209), .C2(new_n212), .ZN(new_n217));
  XOR2_X1   g016(.A(G211gat), .B(G218gat), .Z(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n210), .A2(new_n211), .A3(G204gat), .ZN(new_n221));
  AOI21_X1  g020(.A(G204gat), .B1(new_n210), .B2(new_n211), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n215), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT79), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n203), .A3(new_n215), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n202), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  XOR2_X1   g027(.A(G155gat), .B(G162gat), .Z(new_n229));
  XNOR2_X1  g028(.A(G141gat), .B(G148gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(KEYINPUT2), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT84), .ZN(new_n236));
  OR3_X1    g035(.A1(new_n234), .A2(KEYINPUT84), .A3(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G155gat), .B(G162gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240));
  INV_X1    g039(.A(G162gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT85), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G162gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n240), .B1(new_n245), .B2(G155gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n228), .B(new_n231), .C1(new_n239), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n247), .A2(KEYINPUT87), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT87), .B1(new_n247), .B2(new_n248), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n219), .B1(new_n216), .B2(new_n217), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n225), .A3(new_n218), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT80), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n227), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT88), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT88), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n227), .A2(new_n251), .A3(new_n257), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(G228gat), .A2(G233gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n248), .A3(new_n253), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n228), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n231), .B1(new_n239), .B2(new_n246), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n248), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n227), .A2(new_n254), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n262), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n260), .B2(new_n228), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n259), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G22gat), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n264), .B2(new_n269), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273));
  XNOR2_X1  g072(.A(G78gat), .B(G106gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT31), .B(G50gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NOR4_X1   g076(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n271), .A2(new_n272), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n279), .B2(KEYINPUT89), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n273), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT90), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n227), .A2(new_n254), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NOR3_X1   g085(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  OAI22_X1  g089(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR4_X1   g090(.A1(KEYINPUT71), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  OR2_X1    g096(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  AOI21_X1  g100(.A(G190gat), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n299), .ZN(new_n303));
  NOR2_X1   g102(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n304));
  OAI21_X1  g103(.A(G183gat), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(KEYINPUT69), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT28), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n297), .A2(KEYINPUT27), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT70), .B1(new_n307), .B2(new_n314), .ZN(new_n315));
  AOI211_X1 g114(.A(new_n310), .B(G190gat), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n294), .B(new_n296), .C1(new_n309), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT23), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n321), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  AND2_X1   g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(KEYINPUT23), .B2(new_n319), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n286), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n297), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n286), .A2(KEYINPUT66), .A3(new_n328), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n289), .A2(new_n290), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT67), .B1(new_n338), .B2(new_n321), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n319), .A2(new_n318), .A3(KEYINPUT23), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n326), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n327), .A2(new_n336), .B1(KEYINPUT25), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT29), .B1(new_n317), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT81), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT82), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT83), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n294), .A2(new_n296), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n301), .B(G183gat), .C1(new_n303), .C2(new_n304), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n307), .A2(KEYINPUT69), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n350), .B(new_n332), .C1(new_n300), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n313), .A2(new_n315), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n310), .A2(G190gat), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n352), .A2(new_n310), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n342), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n248), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n346), .ZN(new_n359));
  INV_X1    g158(.A(new_n345), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n285), .A2(new_n348), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n343), .A2(new_n360), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n346), .B1(new_n317), .B2(new_n342), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n284), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n369), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n374), .A3(new_n369), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377));
  XOR2_X1   g176(.A(G113gat), .B(G120gat), .Z(new_n378));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G120gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G113gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT73), .B(G113gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(new_n382), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n379), .B(new_n377), .C1(new_n385), .C2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g185(.A(new_n383), .ZN(new_n387));
  AND2_X1   g186(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n390), .B2(G120gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n381), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n376), .B1(new_n394), .B2(new_n262), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n396), .A3(new_n247), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n379), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n391), .B2(new_n392), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n380), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n267), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n395), .A2(new_n397), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n394), .A2(new_n262), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n267), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n403), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n404), .A2(new_n406), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G1gat), .B(G29gat), .Z(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n412), .B2(new_n413), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n404), .B1(new_n406), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(new_n420), .C1(new_n406), .C2(new_n404), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n373), .A2(new_n375), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT32), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n342), .B(new_n401), .C1(new_n349), .C2(new_n355), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n317), .A2(new_n432), .A3(new_n401), .A4(new_n342), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n356), .A2(new_n394), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT65), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n429), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G71gat), .B(G99gat), .Z(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT33), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n435), .A2(new_n438), .A3(new_n442), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT76), .B1(new_n446), .B2(new_n443), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n447), .B2(new_n439), .ZN(new_n448));
  OR3_X1    g247(.A1(new_n435), .A2(KEYINPUT34), .A3(new_n438), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT34), .B1(new_n435), .B2(new_n437), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n445), .C1(new_n439), .C2(new_n447), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n282), .A2(new_n283), .A3(new_n428), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n264), .A2(new_n269), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G22gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(KEYINPUT89), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n281), .A2(new_n460), .A3(new_n277), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n279), .A2(KEYINPUT89), .A3(new_n276), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n455), .A2(new_n428), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT90), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n464), .A3(KEYINPUT35), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(KEYINPUT90), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n371), .A2(KEYINPUT37), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n372), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n362), .A2(KEYINPUT37), .A3(new_n365), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT38), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n427), .A2(new_n421), .A3(new_n370), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n363), .A2(new_n364), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(new_n285), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n348), .A2(new_n359), .A3(new_n361), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n284), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT38), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n469), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n472), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n395), .A2(new_n402), .A3(new_n397), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n410), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n483), .A2(KEYINPUT39), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n483), .B(KEYINPUT39), .C1(new_n410), .C2(new_n409), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT40), .A4(new_n419), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n419), .B1(new_n483), .B2(KEYINPUT39), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT39), .B1(new_n409), .B2(new_n410), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n410), .B2(new_n482), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n487), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n486), .A2(new_n491), .A3(new_n426), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n373), .A3(new_n375), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n481), .A2(new_n462), .A3(new_n461), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n461), .A2(new_n462), .ZN(new_n495));
  INV_X1    g294(.A(new_n428), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n453), .A2(new_n454), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT77), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT77), .B(KEYINPUT36), .Z(new_n502));
  NAND3_X1  g301(.A1(new_n453), .A2(new_n454), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n494), .A2(new_n497), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n465), .A2(new_n467), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT99), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G155gat), .ZN(new_n509));
  XOR2_X1   g308(.A(G183gat), .B(G211gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G231gat), .ZN(new_n513));
  INV_X1    g312(.A(G233gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(KEYINPUT97), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n519));
  OAI221_X1 g318(.A(new_n517), .B1(G71gat), .B2(G78gat), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n517), .B1(G71gat), .B2(G78gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT98), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT98), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT21), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n516), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G127gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n527), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n533), .A2(KEYINPUT21), .A3(new_n515), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(G1gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT16), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G1gat), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G8gat), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n540), .B(new_n543), .C1(G1gat), .C2(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n545), .B1(new_n533), .B2(KEYINPUT21), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(G127gat), .B1(new_n530), .B2(new_n534), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n536), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(new_n536), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n512), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n549), .A3(new_n511), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT104), .ZN(new_n556));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT41), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT100), .Z(new_n560));
  XOR2_X1   g359(.A(G134gat), .B(G162gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT102), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT103), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G50gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G43gat), .ZN(new_n567));
  INV_X1    g366(.A(G43gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G50gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT15), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OR3_X1    g370(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  NOR3_X1   g373(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G36gat), .ZN(new_n579));
  INV_X1    g378(.A(G29gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT92), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G29gat), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n571), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n570), .A2(KEYINPUT93), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n572), .B1(new_n584), .B2(new_n574), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT15), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n568), .A2(KEYINPUT94), .A3(G50gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n567), .A2(new_n569), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(KEYINPUT94), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n570), .A2(KEYINPUT93), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n586), .A2(new_n587), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  OAI211_X1 g395(.A(KEYINPUT101), .B(KEYINPUT7), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(G85gat), .A3(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n595), .B2(new_n596), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n604), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n558), .B2(new_n557), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n609), .B1(new_n594), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n585), .A2(new_n593), .A3(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n585), .A2(new_n593), .A3(KEYINPUT95), .A4(KEYINPUT17), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n611), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n562), .A2(KEYINPUT102), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n619), .B2(new_n621), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n565), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n619), .A2(new_n621), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n622), .A3(new_n624), .A4(new_n564), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n555), .A2(new_n556), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n556), .B1(new_n555), .B2(new_n629), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n545), .B1(new_n594), .B2(new_n612), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n594), .A2(new_n545), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n585), .A2(new_n593), .B1(new_n542), .B2(new_n544), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n618), .B2(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(KEYINPUT18), .A3(new_n635), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT96), .B1(new_n594), .B2(new_n545), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n542), .A2(new_n544), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n585), .A4(new_n593), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n646), .A3(new_n636), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n635), .B(KEYINPUT13), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n639), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G197gat), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT11), .B(G169gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n639), .A2(new_n655), .A3(new_n642), .A4(new_n649), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n526), .A2(new_n527), .A3(new_n608), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n520), .A2(new_n523), .A3(new_n607), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n606), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n603), .A2(KEYINPUT105), .A3(new_n605), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT106), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT107), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  XOR2_X1   g476(.A(G120gat), .B(G148gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT108), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT10), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n661), .A2(new_n666), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n533), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n668), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n675), .A2(new_n677), .A3(new_n682), .A4(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n681), .B(KEYINPUT109), .Z(new_n689));
  AOI21_X1  g488(.A(new_n669), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n674), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n631), .A2(new_n632), .A3(new_n660), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n506), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n506), .A2(KEYINPUT110), .A3(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n427), .A2(new_n421), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g501(.A1(new_n373), .A2(new_n375), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n698), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n696), .B2(new_n697), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n543), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT42), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(G1325gat));
  INV_X1    g511(.A(new_n698), .ZN(new_n713));
  INV_X1    g512(.A(G15gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(new_n714), .A3(new_n504), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n713), .B2(new_n498), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT111), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n718), .B(new_n714), .C1(new_n713), .C2(new_n498), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(G1326gat));
  NAND2_X1  g519(.A1(new_n698), .A2(new_n495), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT43), .B(G22gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1327gat));
  AND3_X1   g522(.A1(new_n456), .A2(new_n464), .A3(KEYINPUT35), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n505), .A2(new_n467), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n660), .A2(new_n555), .A3(new_n692), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(new_n629), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n581), .A2(new_n583), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n700), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n724), .B2(new_n725), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n465), .A2(KEYINPUT112), .A3(new_n467), .A4(new_n505), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n626), .A2(new_n628), .A3(KEYINPUT113), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT113), .B1(new_n626), .B2(new_n628), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(KEYINPUT44), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n735), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n726), .B2(new_n629), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n699), .B(new_n728), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n733), .B1(new_n731), .B2(new_n743), .ZN(G1328gat));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n579), .A3(new_n704), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n703), .B(new_n728), .C1(new_n741), .C2(new_n742), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n746), .B(new_n747), .C1(new_n579), .C2(new_n748), .ZN(G1329gat));
  NAND2_X1  g548(.A1(new_n741), .A2(new_n742), .ZN(new_n750));
  INV_X1    g549(.A(new_n504), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n750), .A2(G43gat), .A3(new_n751), .A4(new_n727), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n629), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n506), .A2(new_n455), .A3(new_n755), .A4(new_n727), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n756), .A2(new_n568), .B1(KEYINPUT114), .B2(KEYINPUT47), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n752), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n754), .B1(new_n752), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1330gat));
  NOR2_X1   g559(.A1(new_n282), .A2(new_n566), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n750), .A2(new_n727), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n729), .A2(new_n495), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(G50gat), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT48), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n762), .B(new_n766), .C1(G50gat), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1331gat));
  AND2_X1   g567(.A1(new_n735), .A2(new_n736), .ZN(new_n769));
  INV_X1    g568(.A(new_n632), .ZN(new_n770));
  INV_X1    g569(.A(new_n692), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n659), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n770), .A2(new_n630), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n700), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n704), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT49), .B(G64gat), .Z(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(G1333gat));
  NAND4_X1  g579(.A1(new_n769), .A2(G71gat), .A3(new_n751), .A4(new_n773), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n735), .A2(new_n455), .A3(new_n736), .A4(new_n773), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n783));
  INV_X1    g582(.A(G71gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n781), .B(new_n789), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n495), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  INV_X1    g592(.A(new_n555), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n741), .B2(new_n742), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(new_n700), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n555), .A2(new_n659), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n506), .A2(new_n755), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n700), .A2(new_n595), .A3(new_n692), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n797), .A2(new_n595), .B1(new_n804), .B2(new_n805), .ZN(G1336gat));
  AOI21_X1  g605(.A(new_n596), .B1(new_n796), .B2(new_n704), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n703), .A2(new_n771), .A3(G92gat), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n803), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n801), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT52), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n808), .B1(new_n802), .B2(new_n803), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n703), .B(new_n795), .C1(new_n741), .C2(new_n742), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n596), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(G1337gat));
  AND2_X1   g616(.A1(new_n796), .A2(new_n751), .ZN(new_n818));
  INV_X1    g617(.A(G99gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n455), .A2(new_n819), .A3(new_n692), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n818), .A2(new_n819), .B1(new_n804), .B2(new_n820), .ZN(G1338gat));
  INV_X1    g620(.A(G106gat), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n796), .B2(new_n495), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n282), .A2(G106gat), .A3(new_n771), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n810), .B2(new_n801), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n802), .B2(new_n803), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n282), .B(new_n795), .C1(new_n741), .C2(new_n742), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n822), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(G1339gat));
  NOR4_X1   g631(.A1(new_n631), .A2(new_n632), .A3(new_n659), .A4(new_n692), .ZN(new_n833));
  INV_X1    g632(.A(new_n648), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n643), .A2(new_n646), .A3(new_n636), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT116), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n641), .B2(new_n635), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(KEYINPUT116), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n654), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n658), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n684), .A2(new_n669), .A3(new_n685), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n687), .A2(KEYINPUT54), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n682), .B1(new_n690), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(new_n688), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n840), .B(new_n849), .C1(new_n737), .C2(new_n738), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n849), .A2(new_n659), .B1(new_n840), .B2(new_n692), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n739), .B1(new_n851), .B2(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n840), .A2(new_n692), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n847), .A2(new_n688), .A3(new_n848), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n853), .B(KEYINPUT117), .C1(new_n660), .C2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n850), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n833), .B1(new_n857), .B2(new_n794), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n498), .A3(new_n495), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n704), .A2(new_n699), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n660), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(G113gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n384), .B2(new_n862), .ZN(G1340gat));
  NOR2_X1   g663(.A1(new_n861), .A2(new_n771), .ZN(new_n865));
  XOR2_X1   g664(.A(KEYINPUT118), .B(G120gat), .Z(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(G1341gat));
  NOR2_X1   g666(.A1(new_n861), .A2(new_n794), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(new_n532), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n704), .A2(new_n629), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n700), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(G134gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT56), .Z(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n861), .B2(new_n629), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n504), .A2(new_n860), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n282), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n851), .A2(new_n755), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n850), .B1(new_n882), .B2(KEYINPUT120), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n853), .B1(new_n660), .B2(new_n854), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n629), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT121), .B(new_n794), .C1(new_n883), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n833), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n885), .A2(new_n886), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n850), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT121), .B1(new_n893), .B2(new_n794), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n881), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n880), .B1(new_n858), .B2(new_n282), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n879), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n232), .B1(new_n897), .B2(new_n659), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n858), .A2(new_n282), .ZN(new_n899));
  INV_X1    g698(.A(new_n879), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(G141gat), .A3(new_n660), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT58), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(new_n902), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n660), .B(new_n879), .C1(new_n895), .C2(new_n896), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n232), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(G1344gat));
  NAND4_X1  g707(.A1(new_n899), .A2(new_n234), .A3(new_n692), .A4(new_n900), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n884), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n739), .A3(new_n855), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n555), .B1(new_n912), .B2(new_n850), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n881), .B1(new_n913), .B2(new_n833), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n755), .A2(new_n849), .A3(new_n840), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n555), .B1(new_n885), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n495), .B1(new_n916), .B2(new_n833), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n880), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n921));
  AND4_X1   g720(.A1(new_n692), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n234), .B1(new_n897), .B2(new_n692), .ZN(new_n924));
  OAI221_X1 g723(.A(new_n909), .B1(new_n922), .B2(new_n923), .C1(new_n924), .C2(KEYINPUT59), .ZN(G1345gat));
  AND2_X1   g724(.A1(new_n897), .A2(new_n555), .ZN(new_n926));
  INV_X1    g725(.A(G155gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n555), .A2(new_n927), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n926), .A2(new_n927), .B1(new_n901), .B2(new_n928), .ZN(G1346gat));
  NOR3_X1   g728(.A1(new_n873), .A2(new_n245), .A3(new_n751), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n899), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n739), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n897), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n245), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n703), .A2(new_n700), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n859), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n659), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  INV_X1    g739(.A(new_n936), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT123), .B1(new_n941), .B2(new_n498), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n936), .A2(new_n943), .A3(new_n455), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n282), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n858), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n942), .A2(new_n282), .A3(new_n944), .ZN(new_n947));
  OAI211_X1 g746(.A(KEYINPUT124), .B(new_n947), .C1(new_n913), .C2(new_n833), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n660), .A2(new_n289), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n939), .B1(new_n949), .B2(new_n950), .ZN(G1348gat));
  OAI21_X1  g750(.A(new_n290), .B1(new_n937), .B2(new_n771), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n771), .A2(new_n290), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n954), .A2(new_n955), .B1(new_n949), .B2(new_n956), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n946), .A2(new_n555), .A3(new_n948), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G183gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n555), .A2(new_n353), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n937), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g761(.A1(new_n938), .A2(new_n332), .A3(new_n932), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n755), .A3(new_n948), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(G190gat), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n965), .B1(new_n964), .B2(G190gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT61), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n964), .A2(G190gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n972), .B2(new_n966), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n963), .B1(new_n969), .B2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n751), .A2(new_n941), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n899), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n659), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n919), .A2(new_n975), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n660), .A2(new_n207), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  NAND2_X1  g780(.A1(new_n692), .A2(new_n204), .ZN(new_n982));
  OAI21_X1  g781(.A(KEYINPUT62), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  OR3_X1    g782(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n982), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n979), .A2(new_n692), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n204), .ZN(G1353gat));
  INV_X1    g785(.A(G211gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n977), .A2(new_n987), .A3(new_n555), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n979), .A2(new_n555), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  AOI211_X1 g790(.A(new_n991), .B(new_n987), .C1(new_n979), .C2(new_n555), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(G1354gat));
  AOI21_X1  g792(.A(G218gat), .B1(new_n977), .B2(new_n932), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n755), .A2(G218gat), .ZN(new_n995));
  XOR2_X1   g794(.A(new_n995), .B(KEYINPUT127), .Z(new_n996));
  AOI21_X1  g795(.A(new_n994), .B1(new_n979), .B2(new_n996), .ZN(G1355gat));
endmodule


