

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725;

  BUF_X1 U369 ( .A(n627), .Z(n618) );
  NOR2_X1 U370 ( .A1(n725), .A2(n722), .ZN(n352) );
  INV_X2 U371 ( .A(G953), .ZN(n712) );
  XNOR2_X2 U372 ( .A(n358), .B(G113), .ZN(n456) );
  XNOR2_X2 U373 ( .A(n441), .B(n381), .ZN(n709) );
  XOR2_X2 U374 ( .A(KEYINPUT10), .B(n380), .Z(n441) );
  XNOR2_X1 U375 ( .A(n452), .B(n451), .ZN(n597) );
  XOR2_X2 U376 ( .A(G122), .B(G104), .Z(n457) );
  NOR2_X1 U377 ( .A1(n515), .A2(n648), .ZN(n516) );
  XNOR2_X1 U378 ( .A(n492), .B(KEYINPUT40), .ZN(n725) );
  XNOR2_X1 U379 ( .A(n475), .B(n476), .ZN(n722) );
  XNOR2_X1 U380 ( .A(n361), .B(n504), .ZN(n511) );
  NAND2_X1 U381 ( .A1(n509), .A2(n508), .ZN(n518) );
  XNOR2_X1 U382 ( .A(n547), .B(n493), .ZN(n562) );
  XNOR2_X1 U383 ( .A(n565), .B(n499), .ZN(n668) );
  BUF_X1 U384 ( .A(n481), .Z(n547) );
  XNOR2_X1 U385 ( .A(n388), .B(n387), .ZN(n546) );
  NAND2_X1 U386 ( .A1(n597), .A2(n453), .ZN(n360) );
  XNOR2_X1 U387 ( .A(KEYINPUT68), .B(G131), .ZN(n447) );
  XNOR2_X1 U388 ( .A(n522), .B(KEYINPUT73), .ZN(n347) );
  XNOR2_X2 U389 ( .A(n412), .B(n411), .ZN(n508) );
  NOR2_X2 U390 ( .A1(n494), .A2(n667), .ZN(n412) );
  XNOR2_X1 U391 ( .A(n468), .B(n348), .ZN(n497) );
  NAND2_X1 U392 ( .A1(n517), .A2(KEYINPUT47), .ZN(n361) );
  XNOR2_X1 U393 ( .A(n366), .B(KEYINPUT69), .ZN(n365) );
  XNOR2_X1 U394 ( .A(n471), .B(n356), .ZN(n355) );
  INV_X1 U395 ( .A(KEYINPUT112), .ZN(n356) );
  XNOR2_X1 U396 ( .A(n400), .B(KEYINPUT70), .ZN(n494) );
  XNOR2_X1 U397 ( .A(KEYINPUT16), .B(KEYINPUT72), .ZN(n354) );
  XNOR2_X1 U398 ( .A(G119), .B(G110), .ZN(n455) );
  XNOR2_X1 U399 ( .A(n467), .B(n466), .ZN(n630) );
  XNOR2_X1 U400 ( .A(n697), .B(n460), .ZN(n467) );
  NOR2_X1 U401 ( .A1(n569), .A2(n488), .ZN(n489) );
  XNOR2_X1 U402 ( .A(n478), .B(n477), .ZN(n503) );
  XOR2_X1 U403 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n437) );
  NOR2_X1 U404 ( .A1(G953), .A2(G237), .ZN(n446) );
  INV_X1 U405 ( .A(KEYINPUT17), .ZN(n460) );
  XNOR2_X1 U406 ( .A(n363), .B(n362), .ZN(n590) );
  INV_X1 U407 ( .A(KEYINPUT48), .ZN(n362) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n364) );
  XNOR2_X1 U409 ( .A(n528), .B(n469), .ZN(n679) );
  XNOR2_X1 U410 ( .A(n410), .B(G472), .ZN(n481) );
  XNOR2_X1 U411 ( .A(G110), .B(G107), .ZN(n416) );
  XNOR2_X1 U412 ( .A(G104), .B(G101), .ZN(n417) );
  XNOR2_X1 U413 ( .A(n473), .B(n472), .ZN(n677) );
  NAND2_X1 U414 ( .A1(n355), .A2(n680), .ZN(n472) );
  XNOR2_X1 U415 ( .A(n386), .B(n346), .ZN(n387) );
  XNOR2_X1 U416 ( .A(n459), .B(n458), .ZN(n697) );
  XNOR2_X1 U417 ( .A(n353), .B(n455), .ZN(n459) );
  XNOR2_X1 U418 ( .A(n372), .B(n354), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n368), .B(KEYINPUT35), .ZN(n604) );
  NAND2_X1 U420 ( .A1(n370), .A2(n369), .ZN(n368) );
  INV_X1 U421 ( .A(n558), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n371), .B(n350), .ZN(n370) );
  NOR2_X1 U423 ( .A1(n558), .A2(n514), .ZN(n648) );
  INV_X1 U424 ( .A(KEYINPUT105), .ZN(n479) );
  XOR2_X1 U425 ( .A(n385), .B(n384), .Z(n346) );
  AND2_X1 U426 ( .A1(G210), .A2(n470), .ZN(n348) );
  AND2_X1 U427 ( .A1(n550), .A2(n562), .ZN(n349) );
  XOR2_X1 U428 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n350) );
  XOR2_X1 U429 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n351) );
  XNOR2_X2 U430 ( .A(G116), .B(G107), .ZN(n372) );
  NAND2_X1 U431 ( .A1(n355), .A2(n682), .ZN(n683) );
  AND2_X1 U432 ( .A1(n545), .A2(n349), .ZN(n552) );
  XNOR2_X1 U433 ( .A(n544), .B(n357), .ZN(n545) );
  INV_X1 U434 ( .A(KEYINPUT22), .ZN(n357) );
  XNOR2_X2 U435 ( .A(G101), .B(KEYINPUT3), .ZN(n358) );
  NOR2_X4 U436 ( .A1(n359), .A2(n596), .ZN(n627) );
  XNOR2_X2 U437 ( .A(n584), .B(n583), .ZN(n359) );
  NOR2_X1 U438 ( .A1(n663), .A2(n359), .ZN(n693) );
  NAND2_X1 U439 ( .A1(n503), .A2(n502), .ZN(n480) );
  XNOR2_X2 U440 ( .A(n360), .B(n454), .ZN(n478) );
  INV_X1 U441 ( .A(n517), .ZN(n682) );
  AND2_X2 U442 ( .A1(n650), .A2(n652), .ZN(n517) );
  NAND2_X1 U443 ( .A1(n365), .A2(n364), .ZN(n363) );
  NAND2_X1 U444 ( .A1(n347), .A2(n367), .ZN(n366) );
  INV_X1 U445 ( .A(n720), .ZN(n367) );
  NAND2_X1 U446 ( .A1(n557), .A2(n685), .ZN(n371) );
  XNOR2_X1 U447 ( .A(n372), .B(KEYINPUT7), .ZN(n427) );
  XNOR2_X1 U448 ( .A(n506), .B(n505), .ZN(n539) );
  BUF_X1 U449 ( .A(n497), .Z(n528) );
  NAND2_X1 U450 ( .A1(n539), .A2(n538), .ZN(n542) );
  INV_X1 U451 ( .A(KEYINPUT83), .ZN(n504) );
  XNOR2_X1 U452 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U453 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U454 ( .A1(n679), .A2(n678), .ZN(n471) );
  INV_X1 U455 ( .A(KEYINPUT74), .ZN(n583) );
  INV_X1 U456 ( .A(KEYINPUT38), .ZN(n469) );
  BUF_X1 U457 ( .A(n586), .Z(n699) );
  INV_X1 U458 ( .A(KEYINPUT103), .ZN(n477) );
  XNOR2_X1 U459 ( .A(KEYINPUT75), .B(n489), .ZN(n490) );
  INV_X1 U460 ( .A(KEYINPUT60), .ZN(n602) );
  XOR2_X1 U461 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n476) );
  NAND2_X1 U462 ( .A1(n712), .A2(G234), .ZN(n374) );
  XNOR2_X1 U463 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n373) );
  XNOR2_X1 U464 ( .A(n374), .B(n373), .ZN(n425) );
  NAND2_X1 U465 ( .A1(G221), .A2(n425), .ZN(n376) );
  XOR2_X1 U466 ( .A(KEYINPUT78), .B(KEYINPUT24), .Z(n375) );
  XNOR2_X1 U467 ( .A(n376), .B(n375), .ZN(n379) );
  XNOR2_X1 U468 ( .A(G128), .B(KEYINPUT23), .ZN(n377) );
  XNOR2_X1 U469 ( .A(n455), .B(n377), .ZN(n378) );
  XNOR2_X1 U470 ( .A(n379), .B(n378), .ZN(n382) );
  XNOR2_X1 U471 ( .A(G146), .B(G125), .ZN(n462) );
  INV_X1 U472 ( .A(n462), .ZN(n380) );
  XNOR2_X1 U473 ( .A(G140), .B(G137), .ZN(n414) );
  INV_X1 U474 ( .A(n414), .ZN(n381) );
  XNOR2_X1 U475 ( .A(n382), .B(n709), .ZN(n611) );
  NOR2_X1 U476 ( .A1(G902), .A2(n611), .ZN(n388) );
  XNOR2_X1 U477 ( .A(G902), .B(KEYINPUT15), .ZN(n592) );
  NAND2_X1 U478 ( .A1(n592), .A2(G234), .ZN(n383) );
  XNOR2_X1 U479 ( .A(n383), .B(KEYINPUT20), .ZN(n396) );
  NAND2_X1 U480 ( .A1(G217), .A2(n396), .ZN(n386) );
  XOR2_X1 U481 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n385) );
  XNOR2_X1 U482 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n384) );
  NAND2_X1 U483 ( .A1(G234), .A2(G237), .ZN(n389) );
  XNOR2_X1 U484 ( .A(n389), .B(KEYINPUT90), .ZN(n390) );
  XNOR2_X1 U485 ( .A(KEYINPUT14), .B(n390), .ZN(n392) );
  NAND2_X1 U486 ( .A1(n392), .A2(G952), .ZN(n391) );
  XOR2_X1 U487 ( .A(KEYINPUT91), .B(n391), .Z(n691) );
  NOR2_X1 U488 ( .A1(G953), .A2(n691), .ZN(n536) );
  NAND2_X1 U489 ( .A1(n392), .A2(G902), .ZN(n393) );
  XOR2_X1 U490 ( .A(n393), .B(KEYINPUT93), .Z(n533) );
  OR2_X1 U491 ( .A1(n712), .A2(n533), .ZN(n394) );
  NOR2_X1 U492 ( .A1(G900), .A2(n394), .ZN(n395) );
  NOR2_X1 U493 ( .A1(n536), .A2(n395), .ZN(n484) );
  NOR2_X1 U494 ( .A1(n546), .A2(n484), .ZN(n399) );
  NAND2_X1 U495 ( .A1(n396), .A2(G221), .ZN(n398) );
  XOR2_X1 U496 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n397) );
  XNOR2_X1 U497 ( .A(n398), .B(n397), .ZN(n664) );
  NAND2_X1 U498 ( .A1(n399), .A2(n664), .ZN(n400) );
  XOR2_X1 U499 ( .A(G137), .B(KEYINPUT99), .Z(n402) );
  NAND2_X1 U500 ( .A1(n446), .A2(G210), .ZN(n401) );
  XNOR2_X1 U501 ( .A(n402), .B(n401), .ZN(n406) );
  XNOR2_X1 U502 ( .A(G116), .B(G119), .ZN(n404) );
  INV_X1 U503 ( .A(KEYINPUT5), .ZN(n403) );
  XNOR2_X1 U504 ( .A(n456), .B(n407), .ZN(n409) );
  XNOR2_X1 U505 ( .A(n447), .B(G134), .ZN(n408) );
  XNOR2_X2 U506 ( .A(G143), .B(G128), .ZN(n430) );
  XNOR2_X1 U507 ( .A(n430), .B(KEYINPUT4), .ZN(n463) );
  XNOR2_X1 U508 ( .A(n408), .B(n463), .ZN(n710) );
  XNOR2_X1 U509 ( .A(n710), .B(G146), .ZN(n421) );
  XNOR2_X1 U510 ( .A(n409), .B(n421), .ZN(n606) );
  INV_X1 U511 ( .A(G902), .ZN(n453) );
  NAND2_X1 U512 ( .A1(n606), .A2(n453), .ZN(n410) );
  INV_X1 U513 ( .A(n547), .ZN(n667) );
  XOR2_X1 U514 ( .A(KEYINPUT111), .B(KEYINPUT28), .Z(n411) );
  NAND2_X1 U515 ( .A1(n712), .A2(G227), .ZN(n413) );
  XNOR2_X1 U516 ( .A(n413), .B(KEYINPUT79), .ZN(n415) );
  XNOR2_X1 U517 ( .A(n415), .B(n414), .ZN(n419) );
  XNOR2_X1 U518 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U519 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U520 ( .A(n421), .B(n420), .ZN(n622) );
  OR2_X1 U521 ( .A1(n622), .A2(G902), .ZN(n424) );
  INV_X1 U522 ( .A(KEYINPUT71), .ZN(n422) );
  XNOR2_X1 U523 ( .A(n422), .B(G469), .ZN(n423) );
  XNOR2_X2 U524 ( .A(n424), .B(n423), .ZN(n565) );
  XNOR2_X1 U525 ( .A(KEYINPUT110), .B(n565), .ZN(n507) );
  AND2_X1 U526 ( .A1(n508), .A2(n507), .ZN(n474) );
  XOR2_X1 U527 ( .A(KEYINPUT41), .B(KEYINPUT113), .Z(n473) );
  NAND2_X1 U528 ( .A1(G217), .A2(n425), .ZN(n426) );
  XNOR2_X1 U529 ( .A(n427), .B(n426), .ZN(n434) );
  INV_X1 U530 ( .A(G134), .ZN(n428) );
  XNOR2_X1 U531 ( .A(n428), .B(G122), .ZN(n429) );
  XNOR2_X1 U532 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U533 ( .A(KEYINPUT9), .B(KEYINPUT104), .ZN(n431) );
  XNOR2_X1 U534 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U535 ( .A(n434), .B(n433), .ZN(n614) );
  NAND2_X1 U536 ( .A1(n614), .A2(n453), .ZN(n435) );
  XNOR2_X1 U537 ( .A(n435), .B(G478), .ZN(n512) );
  XNOR2_X1 U538 ( .A(n457), .B(KEYINPUT11), .ZN(n439) );
  XNOR2_X1 U539 ( .A(G140), .B(KEYINPUT101), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U542 ( .A1(n441), .A2(n440), .ZN(n445) );
  INV_X1 U543 ( .A(n440), .ZN(n443) );
  INV_X1 U544 ( .A(n441), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X1 U546 ( .A1(n445), .A2(n444), .ZN(n452) );
  NAND2_X1 U547 ( .A1(G214), .A2(n446), .ZN(n448) );
  XNOR2_X1 U548 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U549 ( .A(G113), .B(G143), .ZN(n449) );
  XOR2_X1 U550 ( .A(n450), .B(n449), .Z(n451) );
  XOR2_X1 U551 ( .A(KEYINPUT13), .B(G475), .Z(n454) );
  NOR2_X1 U552 ( .A1(n512), .A2(n478), .ZN(n680) );
  XNOR2_X1 U553 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U554 ( .A1(G224), .A2(n712), .ZN(n461) );
  XNOR2_X1 U555 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U556 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U557 ( .A(n465), .B(KEYINPUT18), .Z(n466) );
  NAND2_X1 U558 ( .A1(n630), .A2(n592), .ZN(n468) );
  OR2_X1 U559 ( .A1(G237), .A2(G902), .ZN(n470) );
  NAND2_X1 U560 ( .A1(G214), .A2(n470), .ZN(n678) );
  NAND2_X1 U561 ( .A1(n474), .A2(n677), .ZN(n475) );
  INV_X1 U562 ( .A(n512), .ZN(n502) );
  XNOR2_X2 U563 ( .A(n480), .B(n479), .ZN(n650) );
  INV_X1 U564 ( .A(n650), .ZN(n496) );
  NAND2_X1 U565 ( .A1(n546), .A2(n664), .ZN(n569) );
  NAND2_X1 U566 ( .A1(n481), .A2(n678), .ZN(n483) );
  XNOR2_X1 U567 ( .A(KEYINPUT30), .B(KEYINPUT109), .ZN(n482) );
  XNOR2_X1 U568 ( .A(n483), .B(n482), .ZN(n487) );
  INV_X1 U569 ( .A(n484), .ZN(n485) );
  AND2_X1 U570 ( .A1(n565), .A2(n485), .ZN(n486) );
  NAND2_X1 U571 ( .A1(n487), .A2(n486), .ZN(n488) );
  INV_X1 U572 ( .A(n490), .ZN(n513) );
  AND2_X1 U573 ( .A1(n513), .A2(n679), .ZN(n491) );
  XOR2_X1 U574 ( .A(n491), .B(KEYINPUT39), .Z(n530) );
  AND2_X1 U575 ( .A1(n496), .A2(n530), .ZN(n492) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT6), .ZN(n493) );
  NOR2_X1 U577 ( .A1(n562), .A2(n494), .ZN(n495) );
  NAND2_X1 U578 ( .A1(n496), .A2(n495), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n497), .A2(n678), .ZN(n506) );
  NOR2_X1 U580 ( .A1(n523), .A2(n506), .ZN(n498) );
  XNOR2_X1 U581 ( .A(KEYINPUT36), .B(n498), .ZN(n500) );
  XNOR2_X1 U582 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n499) );
  INV_X1 U583 ( .A(n668), .ZN(n570) );
  NAND2_X1 U584 ( .A1(n500), .A2(n570), .ZN(n501) );
  XNOR2_X1 U585 ( .A(n501), .B(KEYINPUT115), .ZN(n720) );
  NOR2_X1 U586 ( .A1(n503), .A2(n502), .ZN(n529) );
  INV_X1 U587 ( .A(n529), .ZN(n652) );
  XNOR2_X1 U588 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n505) );
  AND2_X1 U589 ( .A1(n539), .A2(n507), .ZN(n509) );
  NAND2_X1 U590 ( .A1(n518), .A2(KEYINPUT47), .ZN(n510) );
  NAND2_X1 U591 ( .A1(n511), .A2(n510), .ZN(n515) );
  NAND2_X1 U592 ( .A1(n478), .A2(n512), .ZN(n558) );
  NAND2_X1 U593 ( .A1(n528), .A2(n513), .ZN(n514) );
  XNOR2_X1 U594 ( .A(n516), .B(KEYINPUT82), .ZN(n521) );
  XOR2_X1 U595 ( .A(KEYINPUT84), .B(n517), .Z(n576) );
  NOR2_X1 U596 ( .A1(n518), .A2(KEYINPUT47), .ZN(n519) );
  NAND2_X1 U597 ( .A1(n576), .A2(n519), .ZN(n520) );
  NAND2_X1 U598 ( .A1(n521), .A2(n520), .ZN(n522) );
  INV_X1 U599 ( .A(n523), .ZN(n524) );
  NAND2_X1 U600 ( .A1(n524), .A2(n678), .ZN(n525) );
  NOR2_X1 U601 ( .A1(n525), .A2(n570), .ZN(n526) );
  XNOR2_X1 U602 ( .A(n526), .B(KEYINPUT43), .ZN(n527) );
  NOR2_X1 U603 ( .A1(n528), .A2(n527), .ZN(n656) );
  INV_X1 U604 ( .A(n656), .ZN(n531) );
  NAND2_X1 U605 ( .A1(n530), .A2(n529), .ZN(n655) );
  NAND2_X1 U606 ( .A1(n531), .A2(n655), .ZN(n588) );
  INV_X1 U607 ( .A(KEYINPUT2), .ZN(n659) );
  NOR2_X1 U608 ( .A1(n588), .A2(n659), .ZN(n532) );
  AND2_X1 U609 ( .A1(n590), .A2(n532), .ZN(n582) );
  XOR2_X1 U610 ( .A(KEYINPUT92), .B(G898), .Z(n703) );
  NAND2_X1 U611 ( .A1(G953), .A2(n703), .ZN(n698) );
  NOR2_X1 U612 ( .A1(n533), .A2(n698), .ZN(n534) );
  XNOR2_X1 U613 ( .A(n534), .B(KEYINPUT94), .ZN(n535) );
  NOR2_X1 U614 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U615 ( .A(KEYINPUT95), .B(n537), .ZN(n538) );
  INV_X1 U616 ( .A(KEYINPUT88), .ZN(n540) );
  XNOR2_X1 U617 ( .A(n540), .B(KEYINPUT0), .ZN(n541) );
  XNOR2_X2 U618 ( .A(n542), .B(n541), .ZN(n557) );
  AND2_X1 U619 ( .A1(n664), .A2(n680), .ZN(n543) );
  NAND2_X1 U620 ( .A1(n557), .A2(n543), .ZN(n544) );
  NAND2_X1 U621 ( .A1(n545), .A2(n668), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n561), .B(KEYINPUT107), .ZN(n549) );
  NOR2_X1 U623 ( .A1(n546), .A2(n547), .ZN(n548) );
  NAND2_X1 U624 ( .A1(n549), .A2(n548), .ZN(n644) );
  NOR2_X1 U625 ( .A1(n668), .A2(n546), .ZN(n550) );
  INV_X1 U626 ( .A(KEYINPUT32), .ZN(n551) );
  XNOR2_X1 U627 ( .A(n552), .B(n551), .ZN(n723) );
  NAND2_X1 U628 ( .A1(n644), .A2(n723), .ZN(n559) );
  NOR2_X1 U629 ( .A1(n569), .A2(n668), .ZN(n554) );
  INV_X1 U630 ( .A(n562), .ZN(n553) );
  NAND2_X1 U631 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U632 ( .A(KEYINPUT108), .B(KEYINPUT33), .ZN(n555) );
  XNOR2_X1 U633 ( .A(n556), .B(n555), .ZN(n685) );
  NOR2_X2 U634 ( .A1(n559), .A2(n604), .ZN(n560) );
  XNOR2_X1 U635 ( .A(n560), .B(KEYINPUT44), .ZN(n579) );
  INV_X1 U636 ( .A(n561), .ZN(n564) );
  AND2_X1 U637 ( .A1(n562), .A2(n546), .ZN(n563) );
  NAND2_X1 U638 ( .A1(n564), .A2(n563), .ZN(n637) );
  INV_X1 U639 ( .A(n557), .ZN(n572) );
  INV_X1 U640 ( .A(n569), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U642 ( .A1(n572), .A2(n567), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n568), .A2(n667), .ZN(n641) );
  NOR2_X1 U644 ( .A1(n569), .A2(n667), .ZN(n571) );
  NAND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n673) );
  NOR2_X1 U646 ( .A1(n572), .A2(n673), .ZN(n574) );
  XNOR2_X1 U647 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n574), .B(n573), .ZN(n653) );
  NAND2_X1 U649 ( .A1(n641), .A2(n653), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  AND2_X1 U651 ( .A1(n637), .A2(n577), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n581), .B(n580), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n582), .A2(n699), .ZN(n584) );
  INV_X1 U656 ( .A(n592), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT86), .ZN(n591) );
  INV_X1 U659 ( .A(n588), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n711) );
  NOR2_X1 U661 ( .A1(n591), .A2(n711), .ZN(n595) );
  NOR2_X1 U662 ( .A1(n592), .A2(n659), .ZN(n593) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT66), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n627), .A2(G475), .ZN(n599) );
  XOR2_X1 U666 ( .A(n597), .B(KEYINPUT59), .Z(n598) );
  XNOR2_X1 U667 ( .A(n599), .B(n598), .ZN(n601) );
  INV_X1 U668 ( .A(G952), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n600), .A2(G953), .ZN(n633) );
  NAND2_X1 U670 ( .A1(n601), .A2(n633), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(n602), .ZN(G60) );
  XOR2_X1 U672 ( .A(G122), .B(n604), .Z(G24) );
  NAND2_X1 U673 ( .A1(n627), .A2(G472), .ZN(n608) );
  XOR2_X1 U674 ( .A(KEYINPUT89), .B(KEYINPUT62), .Z(n605) );
  XNOR2_X1 U675 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U676 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n609), .A2(n633), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n610), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U679 ( .A1(n618), .A2(G217), .ZN(n612) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n613) );
  INV_X1 U681 ( .A(n633), .ZN(n625) );
  NOR2_X1 U682 ( .A1(n613), .A2(n625), .ZN(G66) );
  NAND2_X1 U683 ( .A1(n618), .A2(G478), .ZN(n616) );
  XNOR2_X1 U684 ( .A(n614), .B(KEYINPUT123), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X1 U686 ( .A1(n617), .A2(n625), .ZN(G63) );
  NAND2_X1 U687 ( .A1(n618), .A2(G469), .ZN(n624) );
  XNOR2_X1 U688 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n620) );
  XNOR2_X1 U689 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(n626) );
  NOR2_X1 U693 ( .A1(n626), .A2(n625), .ZN(G54) );
  NAND2_X1 U694 ( .A1(n627), .A2(G210), .ZN(n632) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT55), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U698 ( .A(n632), .B(n631), .ZN(n634) );
  NAND2_X1 U699 ( .A1(n634), .A2(n633), .ZN(n636) );
  XOR2_X1 U700 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n635) );
  XNOR2_X1 U701 ( .A(n636), .B(n635), .ZN(G51) );
  XNOR2_X1 U702 ( .A(G101), .B(n637), .ZN(G3) );
  NOR2_X1 U703 ( .A1(n650), .A2(n641), .ZN(n638) );
  XOR2_X1 U704 ( .A(G104), .B(n638), .Z(G6) );
  XOR2_X1 U705 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  XNOR2_X1 U706 ( .A(G107), .B(KEYINPUT116), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(n643) );
  NOR2_X1 U708 ( .A1(n652), .A2(n641), .ZN(n642) );
  XOR2_X1 U709 ( .A(n643), .B(n642), .Z(G9) );
  XNOR2_X1 U710 ( .A(n644), .B(G110), .ZN(G12) );
  NOR2_X1 U711 ( .A1(n652), .A2(n518), .ZN(n646) );
  XNOR2_X1 U712 ( .A(KEYINPUT117), .B(KEYINPUT29), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U714 ( .A(G128), .B(n647), .Z(G30) );
  XOR2_X1 U715 ( .A(G143), .B(n648), .Z(G45) );
  NOR2_X1 U716 ( .A1(n650), .A2(n518), .ZN(n649) );
  XOR2_X1 U717 ( .A(G146), .B(n649), .Z(G48) );
  NOR2_X1 U718 ( .A1(n653), .A2(n650), .ZN(n651) );
  XOR2_X1 U719 ( .A(G113), .B(n651), .Z(G15) );
  NOR2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U721 ( .A(G116), .B(n654), .Z(G18) );
  XNOR2_X1 U722 ( .A(G134), .B(n655), .ZN(G36) );
  XOR2_X1 U723 ( .A(G140), .B(n656), .Z(n657) );
  XNOR2_X1 U724 ( .A(KEYINPUT118), .B(n657), .ZN(G42) );
  AND2_X1 U725 ( .A1(n677), .A2(n685), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n658), .A2(G953), .ZN(n695) );
  NAND2_X1 U727 ( .A1(n711), .A2(n659), .ZN(n660) );
  XOR2_X1 U728 ( .A(n660), .B(KEYINPUT85), .Z(n662) );
  OR2_X1 U729 ( .A1(n699), .A2(KEYINPUT2), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n664), .A2(n546), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n665), .B(KEYINPUT49), .ZN(n666) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n569), .A2(n668), .ZN(n669) );
  XOR2_X1 U735 ( .A(KEYINPUT50), .B(n669), .Z(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT119), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n675), .Z(n676) );
  NAND2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n688) );
  OR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n684) );
  NAND2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n689), .Z(n690) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(n696), .Z(G75) );
  NAND2_X1 U751 ( .A1(n698), .A2(n697), .ZN(n708) );
  NAND2_X1 U752 ( .A1(n699), .A2(n712), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n700), .B(KEYINPUT125), .ZN(n706) );
  NAND2_X1 U754 ( .A1(G953), .A2(G224), .ZN(n701) );
  XOR2_X1 U755 ( .A(KEYINPUT61), .B(n701), .Z(n702) );
  NOR2_X1 U756 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U757 ( .A(KEYINPUT124), .B(n704), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(G69) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(n715) );
  XNOR2_X1 U761 ( .A(n711), .B(n715), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n714), .B(KEYINPUT126), .ZN(n719) );
  XNOR2_X1 U764 ( .A(n715), .B(G227), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n716), .A2(G900), .ZN(n717) );
  NAND2_X1 U766 ( .A1(G953), .A2(n717), .ZN(n718) );
  NAND2_X1 U767 ( .A1(n719), .A2(n718), .ZN(G72) );
  XNOR2_X1 U768 ( .A(G125), .B(n720), .ZN(n721) );
  XNOR2_X1 U769 ( .A(n721), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U770 ( .A(n722), .B(G137), .Z(G39) );
  XOR2_X1 U771 ( .A(G119), .B(n723), .Z(n724) );
  XNOR2_X1 U772 ( .A(KEYINPUT127), .B(n724), .ZN(G21) );
  XOR2_X1 U773 ( .A(G131), .B(n725), .Z(G33) );
endmodule

