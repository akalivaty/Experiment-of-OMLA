//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(G1gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(G1gat), .ZN(new_n209));
  OAI21_X1  g008(.A(G8gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n211), .B(new_n212), .C1(G1gat), .C2(new_n205), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT89), .B(G36gat), .Z(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G29gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT88), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n219), .B(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT88), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT15), .B(new_n216), .C1(new_n222), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G50gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT90), .B1(new_n227), .B2(G43gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT15), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(new_n216), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(new_n224), .A3(new_n218), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n226), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n226), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n215), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n226), .A2(new_n231), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n210), .B2(new_n213), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n202), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n233), .A2(new_n234), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n237), .B1(new_n244), .B2(new_n215), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(KEYINPUT18), .A3(new_n240), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n215), .A2(new_n236), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n238), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n240), .B(KEYINPUT13), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n242), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT11), .B(G169gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G197gat), .ZN(new_n254));
  XOR2_X1   g053(.A(G113gat), .B(G141gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT12), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n242), .A2(new_n246), .A3(new_n257), .A4(new_n251), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT35), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(G183gat), .B2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n280), .A2(G169gat), .A3(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT25), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n286), .B(new_n270), .C1(new_n272), .C2(new_n274), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n276), .A2(new_n281), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT66), .B1(new_n282), .B2(new_n284), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290));
  OAI211_X1 g089(.A(G183gat), .B(G190gat), .C1(new_n290), .C2(KEYINPUT24), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n273), .A2(KEYINPUT67), .A3(new_n271), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n270), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(new_n283), .C1(new_n279), .C2(new_n280), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n289), .A2(new_n293), .A3(new_n295), .A4(new_n281), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT25), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n279), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(KEYINPUT26), .B2(new_n279), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n284), .A2(KEYINPUT70), .B1(new_n279), .B2(KEYINPUT26), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n268), .A2(KEYINPUT27), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n304), .B1(new_n306), .B2(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n269), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n303), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(new_n303), .C1(new_n308), .C2(new_n310), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n305), .A2(new_n307), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n269), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n298), .B1(new_n302), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n319), .A2(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G127gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n321), .A2(G127gat), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT71), .B(G127gat), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT72), .B(new_n322), .C1(new_n326), .C2(new_n321), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n329), .A2(KEYINPUT71), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(KEYINPUT71), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n328), .B(G134gat), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n327), .A2(KEYINPUT73), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT73), .B1(new_n327), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n325), .B1(new_n335), .B2(new_n320), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT75), .B1(new_n318), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n302), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n288), .A2(new_n297), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n322), .A2(KEYINPUT72), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT71), .B(G127gat), .Z(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(G134gat), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n326), .A2(KEYINPUT72), .A3(new_n321), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n327), .A2(KEYINPUT73), .A3(new_n332), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n320), .ZN(new_n349));
  INV_X1    g148(.A(new_n325), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n340), .A2(new_n341), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT74), .B1(new_n340), .B2(new_n351), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n336), .A2(new_n355), .A3(new_n338), .A4(new_n339), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n359), .B(KEYINPUT64), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n267), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n337), .A2(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT32), .B1(new_n366), .B2(new_n360), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n361), .A2(KEYINPUT34), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT77), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AND4_X1   g168(.A1(KEYINPUT77), .A2(new_n353), .A3(new_n357), .A4(new_n368), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n357), .A3(new_n368), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n368), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n367), .A2(new_n378), .A3(new_n374), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n365), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT31), .B(G50gat), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT78), .B(G211gat), .Z(new_n384));
  AOI21_X1  g183(.A(KEYINPUT22), .B1(new_n384), .B2(G218gat), .ZN(new_n385));
  XOR2_X1   g184(.A(G197gat), .B(G204gat), .Z(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n388));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  XNOR2_X1  g189(.A(G155gat), .B(G162gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G141gat), .B(G148gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(KEYINPUT2), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  INV_X1    g194(.A(G162gat), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT2), .B1(new_n396), .B2(KEYINPUT82), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n390), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n388), .B(new_n389), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n403), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n400), .B1(new_n410), .B2(new_n401), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n406), .B(KEYINPUT85), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n387), .B2(new_n389), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n387), .B2(new_n389), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n401), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n399), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n405), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n383), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G78gat), .B(G106gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G22gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n413), .ZN(new_n424));
  INV_X1    g223(.A(new_n383), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n424), .B(new_n425), .C1(new_n411), .C2(new_n408), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n420), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n422), .B1(new_n420), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n318), .B2(KEYINPUT29), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n390), .C1(new_n318), .C2(new_n430), .ZN(new_n432));
  INV_X1    g231(.A(new_n430), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n340), .B2(new_n403), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n318), .A2(new_n430), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n409), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G8gat), .B(G36gat), .Z(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G64gat), .ZN(new_n439));
  INV_X1    g238(.A(G92gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT81), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n441), .B1(new_n432), .B2(new_n436), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT30), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(KEYINPUT30), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n441), .B(KEYINPUT80), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n436), .A3(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n378), .A2(new_n374), .A3(new_n379), .ZN(new_n454));
  INV_X1    g253(.A(new_n367), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n364), .A3(new_n380), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n382), .A2(new_n429), .A3(new_n453), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n399), .A2(KEYINPUT3), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n351), .A2(new_n402), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n349), .A2(new_n400), .A3(new_n350), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT4), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n349), .A2(new_n467), .A3(new_n400), .A4(new_n350), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n465), .B2(new_n468), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n460), .B(new_n463), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n464), .A4(new_n461), .ZN(new_n472));
  INV_X1    g271(.A(new_n464), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n400), .B1(new_n349), .B2(new_n350), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT5), .A4(new_n468), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT0), .B(G57gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(G85gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  NAND3_X1  g279(.A1(new_n471), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n471), .B2(new_n476), .ZN(new_n484));
  MUX2_X1   g283(.A(new_n483), .B(new_n482), .S(new_n484), .Z(new_n485));
  OAI21_X1  g284(.A(new_n263), .B1(new_n458), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n456), .A2(new_n364), .A3(new_n380), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n364), .B1(new_n456), .B2(new_n380), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT84), .B1(new_n481), .B2(new_n482), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n484), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n481), .A2(KEYINPUT84), .A3(new_n482), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(KEYINPUT6), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n263), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n489), .A2(new_n496), .A3(new_n429), .A4(new_n453), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n487), .B2(new_n488), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n382), .A2(KEYINPUT36), .A3(new_n457), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n437), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT37), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n441), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n447), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n450), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n507), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n504), .A2(new_n513), .A3(new_n505), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n485), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n462), .ZN(new_n518));
  OR3_X1    g317(.A1(new_n473), .A2(new_n462), .A3(new_n474), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(KEYINPUT39), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT39), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n521), .A3(new_n462), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n480), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT40), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n520), .A2(KEYINPUT40), .A3(new_n480), .A4(new_n522), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n452), .A3(new_n526), .A4(new_n492), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n516), .A2(new_n429), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n429), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n493), .A2(new_n492), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n495), .B1(new_n530), .B2(new_n490), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n532), .B2(new_n452), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n502), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n262), .B1(new_n498), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT9), .ZN(new_n537));
  INV_X1    g336(.A(G71gat), .ZN(new_n538));
  INV_X1    g337(.A(G78gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(KEYINPUT94), .B(new_n540), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n536), .B(KEYINPUT92), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  OAI221_X1 g349(.A(new_n549), .B1(new_n550), .B2(new_n541), .C1(new_n538), .C2(new_n539), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n214), .B1(new_n553), .B2(KEYINPUT21), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(new_n268), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n553), .A2(KEYINPUT21), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n559), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G211gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n560), .A2(new_n568), .A3(new_n561), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G190gat), .B(G218gat), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT100), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n576), .B1(new_n577), .B2(new_n440), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n577), .B2(new_n440), .ZN(new_n580));
  NAND3_X1  g379(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT98), .ZN(new_n583));
  XOR2_X1   g382(.A(G99gat), .B(G106gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n582), .A2(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(KEYINPUT98), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(new_n236), .C1(new_n592), .C2(KEYINPUT17), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n236), .A2(new_n232), .ZN(new_n594));
  INV_X1    g393(.A(new_n234), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT99), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n593), .B1(new_n596), .B2(new_n591), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n574), .A2(KEYINPUT100), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n599));
  AND4_X1   g398(.A1(new_n321), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n590), .B1(new_n243), .B2(KEYINPUT99), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(new_n593), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n321), .B1(new_n603), .B2(new_n598), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n575), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(G134gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n575), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n321), .A3(new_n598), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT97), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G162gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n614), .A3(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n552), .A2(new_n590), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n548), .A2(new_n586), .A3(new_n551), .A4(new_n589), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G230gat), .ZN(new_n622));
  INV_X1    g421(.A(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n627), .A3(new_n620), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n553), .A2(new_n591), .A3(KEYINPUT10), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(new_n278), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(G204gat), .Z(new_n633));
  OR3_X1    g432(.A1(new_n626), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n626), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n572), .A2(new_n618), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n535), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n531), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT101), .B(G1gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1324gat));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n453), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n206), .A2(new_n212), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n645), .A2(KEYINPUT42), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(KEYINPUT42), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n646), .B(new_n647), .C1(new_n212), .C2(new_n642), .ZN(G1325gat));
  INV_X1    g447(.A(G15gat), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n638), .A2(new_n649), .A3(new_n502), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n535), .A2(new_n489), .A3(new_n637), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n649), .B2(new_n651), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n638), .A2(new_n429), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n570), .A2(new_n571), .ZN(new_n656));
  INV_X1    g455(.A(new_n617), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n614), .B1(new_n605), .B2(new_n610), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n656), .A2(new_n659), .A3(new_n636), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n535), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n532), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(G29gat), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n662), .A2(KEYINPUT102), .A3(G29gat), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n502), .A2(new_n528), .A3(new_n533), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n486), .A2(new_n497), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n618), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT44), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT104), .B1(new_n616), .B2(new_n617), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(KEYINPUT44), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n669), .B2(new_n670), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT105), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n534), .A2(new_n486), .A3(new_n497), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n681), .A3(new_n677), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n672), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n261), .B(KEYINPUT103), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n656), .A2(new_n636), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n531), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n668), .A2(new_n688), .A3(new_n689), .ZN(G1328gat));
  NAND2_X1  g489(.A1(new_n535), .A2(new_n660), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(new_n217), .A3(new_n453), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n217), .B1(new_n687), .B2(new_n453), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1329gat));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n697));
  INV_X1    g496(.A(new_n489), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n691), .A2(G43gat), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n687), .A2(new_n502), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n697), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1330gat));
  OAI21_X1  g503(.A(G50gat), .B1(new_n687), .B2(new_n429), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n429), .B1(new_n661), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n707), .B(new_n227), .C1(new_n706), .C2(new_n661), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g509(.A1(new_n656), .A2(new_n659), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n498), .B2(new_n534), .ZN(new_n712));
  INV_X1    g511(.A(new_n636), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n685), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n532), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g517(.A(new_n453), .B(new_n715), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n719));
  OR2_X1    g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n724), .A3(new_n722), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1333gat));
  NOR3_X1   g527(.A1(new_n715), .A2(new_n538), .A3(new_n502), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n716), .A2(new_n489), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n538), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n429), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n539), .ZN(G1335gat));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(KEYINPUT51), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n656), .A2(new_n685), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n680), .A2(new_n618), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(KEYINPUT51), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n636), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n532), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n683), .A2(new_n572), .A3(new_n714), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n532), .A2(G85gat), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(G1336gat));
  OAI21_X1  g546(.A(new_n440), .B1(new_n741), .B2(new_n453), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(G92gat), .A3(new_n452), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1337gat));
  OR3_X1    g551(.A1(new_n741), .A2(G99gat), .A3(new_n698), .ZN(new_n753));
  INV_X1    g552(.A(new_n502), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G99gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(new_n756), .A3(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1338gat));
  NAND4_X1  g560(.A1(new_n683), .A2(new_n529), .A3(new_n572), .A4(new_n714), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n429), .A2(G106gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n659), .B1(new_n498), .B2(new_n534), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n766), .A2(new_n737), .B1(new_n735), .B2(KEYINPUT51), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n738), .A2(new_n739), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n636), .B(new_n765), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n740), .A2(KEYINPUT112), .A3(new_n636), .A4(new_n765), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n763), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n774), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT113), .B1(new_n774), .B2(KEYINPUT53), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n770), .B1(new_n775), .B2(new_n776), .ZN(G1339gat));
  NOR2_X1   g576(.A1(new_n698), .A2(new_n529), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n245), .B2(new_n240), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n238), .A2(new_n247), .A3(new_n249), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n239), .A2(KEYINPUT115), .A3(new_n241), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n256), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n260), .A3(new_n636), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n628), .A2(new_n629), .A3(new_n624), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n630), .B2(KEYINPUT114), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n628), .A2(new_n629), .A3(new_n788), .A4(new_n624), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n633), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n630), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n634), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n785), .B1(new_n684), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n676), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n260), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n674), .B2(new_n675), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n656), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n711), .A2(new_n636), .A3(new_n685), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n532), .B(new_n778), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n452), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT116), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n806), .B2(new_n452), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n262), .ZN(new_n812));
  INV_X1    g611(.A(new_n807), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n813), .A2(G113gat), .A3(new_n684), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT117), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n811), .B2(new_n713), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n813), .A2(G120gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n713), .B2(new_n821), .ZN(G1341gat));
  OAI21_X1  g621(.A(new_n344), .B1(new_n813), .B2(new_n572), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n656), .A2(new_n326), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n811), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT118), .ZN(G1342gat));
  OAI21_X1  g625(.A(G134gat), .B1(new_n811), .B2(new_n659), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n618), .A2(new_n453), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n806), .A2(G134gat), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT56), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n830), .ZN(G1343gat));
  NAND4_X1  g630(.A1(new_n796), .A2(new_n261), .A3(new_n634), .A4(new_n797), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n785), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n784), .A2(new_n636), .A3(KEYINPUT119), .A4(new_n260), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n659), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n673), .B1(new_n657), .B2(new_n658), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n616), .A2(KEYINPUT104), .A3(new_n617), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n838), .A2(KEYINPUT120), .B1(new_n841), .B2(new_n802), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n835), .A2(new_n836), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n618), .B1(new_n843), .B2(new_n832), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n656), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n529), .C1(new_n847), .C2(new_n805), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n803), .B1(new_n844), .B2(new_n845), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n572), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n805), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n529), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n529), .B1(new_n804), .B2(new_n805), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n850), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n754), .A2(new_n531), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n453), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n261), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G141gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n857), .A2(G141gat), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n261), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT122), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n860), .A2(new_n685), .A3(new_n863), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n871), .A2(G141gat), .B1(new_n261), .B2(new_n866), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(new_n869), .ZN(G1344gat));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n860), .A2(new_n863), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n874), .B(G148gat), .C1(new_n875), .C2(new_n713), .ZN(new_n876));
  XOR2_X1   g675(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n877));
  NAND2_X1  g676(.A1(new_n637), .A2(new_n262), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n802), .A2(new_n618), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n572), .B1(new_n844), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n529), .A2(new_n881), .B1(new_n857), .B2(KEYINPUT57), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(new_n636), .A3(new_n863), .ZN(new_n883));
  INV_X1    g682(.A(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n857), .A2(new_n862), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n884), .A3(new_n636), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1345gat));
  AOI21_X1  g688(.A(G155gat), .B1(new_n887), .B2(new_n656), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n572), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(G155gat), .ZN(G1346gat));
  XOR2_X1   g691(.A(KEYINPUT82), .B(G162gat), .Z(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n875), .B2(new_n676), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n804), .A2(new_n805), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n828), .A2(new_n893), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n895), .A2(new_n529), .A3(new_n861), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n532), .A2(new_n453), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n778), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT124), .Z(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n277), .A3(new_n685), .ZN(new_n902));
  OAI21_X1  g701(.A(G169gat), .B1(new_n900), .B2(new_n262), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1348gat));
  NOR3_X1   g703(.A1(new_n900), .A2(new_n278), .A3(new_n713), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n636), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n278), .ZN(G1349gat));
  OAI21_X1  g706(.A(new_n268), .B1(new_n900), .B2(new_n572), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n900), .A2(new_n572), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n315), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n269), .A3(new_n841), .ZN(new_n912));
  OAI21_X1  g711(.A(G190gat), .B1(new_n900), .B2(new_n659), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT61), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1351gat));
  NAND2_X1  g714(.A1(new_n502), .A2(new_n899), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n882), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n262), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n529), .A3(new_n917), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(G197gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n684), .B2(new_n921), .ZN(G1352gat));
  NOR3_X1   g721(.A1(new_n920), .A2(G204gat), .A3(new_n713), .ZN(new_n923));
  XNOR2_X1  g722(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n882), .A2(new_n636), .A3(new_n917), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G204gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1353gat));
  OAI21_X1  g727(.A(G211gat), .B1(new_n918), .B2(new_n572), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT63), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT63), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n920), .A2(new_n384), .A3(new_n572), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT126), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(G1354gat));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n618), .B1(new_n918), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT127), .B1(new_n882), .B2(new_n917), .ZN(new_n937));
  OAI21_X1  g736(.A(G218gat), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n676), .A2(G218gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n920), .B2(new_n939), .ZN(G1355gat));
endmodule


