//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT80), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(new_n211), .C1(new_n212), .C2(KEYINPUT2), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(KEYINPUT2), .B2(new_n211), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n212), .A2(KEYINPUT74), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n212), .A2(KEYINPUT74), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT75), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n212), .B(KEYINPUT74), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n215), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n214), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT29), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(G211gat), .ZN(new_n227));
  INV_X1    g026(.A(G218gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n226), .B1(KEYINPUT22), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G211gat), .B(G218gat), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT81), .B1(new_n225), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G228gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n218), .A2(KEYINPUT75), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n221), .B1(new_n220), .B2(new_n215), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n224), .B(new_n213), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n232), .B1(new_n240), .B2(new_n235), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n233), .B(new_n234), .C1(new_n237), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n234), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n241), .A2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G22gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n242), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n242), .B2(new_n246), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n205), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n246), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(KEYINPUT82), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n242), .B(new_n246), .C1(KEYINPUT82), .C2(new_n247), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n204), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  INV_X1    g056(.A(G120gat), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n257), .B2(new_n258), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n223), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n262), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT77), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n262), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n223), .B2(new_n224), .ZN(new_n272));
  INV_X1    g071(.A(new_n240), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n213), .B1(new_n238), .B2(new_n239), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n262), .B1(new_n276), .B2(KEYINPUT3), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT76), .B1(new_n277), .B2(new_n240), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n267), .B(new_n270), .C1(new_n275), .C2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n271), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n263), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n280), .B1(new_n283), .B2(new_n269), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n266), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n274), .B1(new_n272), .B2(new_n273), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n277), .A2(KEYINPUT76), .A3(new_n240), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n288), .B2(new_n270), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n291));
  XOR2_X1   g090(.A(G1gat), .B(G29gat), .Z(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G57gat), .B(G85gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n281), .B2(new_n289), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT79), .A3(new_n291), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302));
  INV_X1    g101(.A(new_n284), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n288), .A2(KEYINPUT5), .A3(new_n270), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(KEYINPUT6), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n296), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n298), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT73), .ZN(new_n313));
  XOR2_X1   g112(.A(G64gat), .B(G92gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n232), .ZN(new_n316));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT65), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT24), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT66), .B(G183gat), .Z(new_n325));
  OAI21_X1  g124(.A(new_n324), .B1(G190gat), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT64), .ZN(new_n328));
  INV_X1    g127(.A(new_n319), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n321), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n326), .A2(KEYINPUT25), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n322), .A2(new_n331), .B1(new_n338), .B2(KEYINPUT25), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n325), .A2(KEYINPUT27), .ZN(new_n340));
  OR2_X1    g139(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n341), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n333), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n342), .A2(new_n343), .B1(new_n348), .B2(KEYINPUT28), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n329), .A2(KEYINPUT26), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n328), .B(new_n350), .C1(new_n320), .C2(KEYINPUT26), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n323), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n351), .B2(new_n323), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n339), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n318), .B1(new_n356), .B2(new_n235), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(new_n323), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT68), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n353), .A3(new_n349), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n317), .B1(new_n360), .B2(new_n339), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n316), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n318), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n360), .B2(new_n339), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n363), .B(new_n232), .C1(new_n364), .C2(new_n318), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(KEYINPUT72), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT72), .B1(new_n362), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n315), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n365), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(new_n315), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n311), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n371), .A2(KEYINPUT30), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n256), .B1(new_n310), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT36), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n378));
  INV_X1    g177(.A(G227gat), .ZN(new_n379));
  INV_X1    g178(.A(G233gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n339), .B(new_n262), .C1(new_n354), .C2(new_n355), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n262), .B1(new_n360), .B2(new_n339), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G15gat), .B(G43gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT33), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(KEYINPUT32), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT69), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n356), .A2(new_n271), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n382), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n395), .B2(new_n381), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n390), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n385), .A2(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n388), .B1(new_n385), .B2(KEYINPUT32), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n392), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n381), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n402), .A3(new_n382), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n405), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n378), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n398), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n400), .A2(new_n399), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n411), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n401), .A2(KEYINPUT71), .A3(new_n409), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n377), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n391), .A2(KEYINPUT69), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n397), .B1(new_n396), .B2(new_n390), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n412), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n408), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n401), .A2(new_n409), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n377), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT83), .B1(new_n376), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n422), .A3(new_n378), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n415), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n423), .B1(new_n428), .B2(new_n377), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n304), .A2(new_n305), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n299), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n301), .B2(new_n307), .ZN(new_n433));
  INV_X1    g232(.A(new_n374), .ZN(new_n434));
  INV_X1    g233(.A(new_n368), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n366), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n371), .B1(new_n436), .B2(new_n315), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n437), .B2(new_n311), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n433), .A2(new_n438), .A3(new_n298), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n429), .B(new_n430), .C1(new_n439), .C2(new_n256), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT6), .B1(new_n431), .B2(new_n299), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n297), .B1(new_n441), .B2(new_n432), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n435), .B2(new_n366), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n362), .A2(new_n444), .A3(new_n365), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n315), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n447), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n443), .B1(new_n370), .B2(KEYINPUT37), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n371), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT39), .ZN(new_n453));
  INV_X1    g252(.A(new_n283), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n270), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n288), .B2(new_n270), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n267), .B1(new_n275), .B2(new_n278), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n453), .A3(new_n269), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n458), .A3(new_n299), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n296), .A2(new_n290), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n459), .A2(new_n460), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n462), .C1(new_n373), .C2(new_n374), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n452), .A2(new_n463), .A3(new_n256), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n426), .A2(new_n440), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n308), .A2(new_n309), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n421), .A2(new_n256), .A3(new_n422), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n297), .A4(new_n375), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT35), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n438), .A2(new_n442), .A3(KEYINPUT35), .ZN(new_n470));
  INV_X1    g269(.A(new_n256), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n427), .B2(new_n415), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  XNOR2_X1  g275(.A(G71gat), .B(G78gat), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n478));
  INV_X1    g277(.A(G57gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G64gat), .ZN(new_n480));
  INV_X1    g279(.A(G64gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G57gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n476), .B(new_n477), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n482), .ZN(new_n486));
  INV_X1    g285(.A(new_n478), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT89), .B1(new_n488), .B2(KEYINPUT88), .ZN(new_n489));
  INV_X1    g288(.A(new_n477), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n488), .B2(KEYINPUT89), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT21), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G231gat), .A2(G233gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(G127gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT16), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(G1gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G1gat), .B2(new_n498), .ZN(new_n501));
  INV_X1    g300(.A(G8gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n493), .B2(new_n492), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n497), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(new_n206), .ZN(new_n507));
  XOR2_X1   g306(.A(G183gat), .B(G211gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n505), .A2(new_n510), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(G29gat), .ZN(new_n518));
  INV_X1    g317(.A(G36gat), .ZN(new_n519));
  OAI22_X1  g318(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT15), .A3(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n521), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(KEYINPUT15), .B2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n517), .A2(new_n525), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n516), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n522), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT17), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT91), .A2(G92gat), .ZN(new_n531));
  INV_X1    g330(.A(G85gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(KEYINPUT91), .A2(G92gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G99gat), .ZN(new_n535));
  INV_X1    g334(.A(G106gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT8), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(KEYINPUT90), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n534), .A2(new_n537), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G99gat), .B(G106gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(KEYINPUT92), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n544), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(new_n543), .A3(new_n537), .A4(new_n534), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n530), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n545), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n529), .ZN(new_n553));
  NAND3_X1  g352(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G190gat), .B(G218gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G134gat), .B(G162gat), .Z(new_n558));
  AOI21_X1  g357(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT93), .Z(new_n561));
  OR2_X1    g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(KEYINPUT93), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n514), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n530), .A2(new_n503), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT87), .Z(new_n569));
  INV_X1    g368(.A(new_n503), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n529), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n503), .B(new_n529), .Z(new_n576));
  XOR2_X1   g375(.A(new_n569), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT85), .B(G197gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT11), .B(G169gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT12), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n579), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n492), .A2(new_n550), .A3(new_n545), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(KEYINPUT10), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT88), .B1(new_n593), .B2(new_n478), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT89), .B1(new_n593), .B2(new_n478), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n476), .A2(new_n594), .B1(new_n595), .B2(new_n477), .ZN(new_n596));
  INV_X1    g395(.A(new_n485), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n546), .A2(new_n548), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n592), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n546), .A2(new_n548), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n492), .A2(new_n601), .A3(KEYINPUT94), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n590), .B(new_n591), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n552), .A2(KEYINPUT10), .A3(new_n598), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n589), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n590), .B1(new_n600), .B2(new_n602), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n589), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G120gat), .B(G148gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n587), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n603), .A2(new_n604), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n588), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n589), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n611), .B1(new_n615), .B2(KEYINPUT96), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(KEYINPUT96), .B2(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n614), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n620), .B1(new_n619), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n566), .A2(new_n586), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n475), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n310), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT100), .B(G1gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1324gat));
  INV_X1    g431(.A(new_n628), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G8gat), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n633), .A2(new_n375), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n502), .B1(new_n628), .B2(new_n438), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT42), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(KEYINPUT42), .B2(new_n636), .ZN(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n633), .B2(new_n429), .ZN(new_n640));
  INV_X1    g439(.A(G15gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n628), .A2(new_n641), .A3(new_n428), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n471), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT43), .B(G22gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  INV_X1    g445(.A(new_n464), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n429), .B1(new_n439), .B2(new_n256), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(KEYINPUT83), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(new_n440), .B1(new_n469), .B2(new_n473), .ZN(new_n650));
  INV_X1    g449(.A(new_n565), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n626), .ZN(new_n653));
  INV_X1    g452(.A(new_n586), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n653), .A2(new_n654), .A3(new_n513), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n518), .A3(new_n629), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT44), .B1(new_n650), .B2(new_n651), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n429), .B(new_n464), .C1(new_n439), .C2(new_n256), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n474), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n474), .A2(new_n661), .A3(new_n660), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n565), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n655), .ZN(new_n668));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668), .B2(new_n310), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(new_n669), .ZN(G1328gat));
  NAND3_X1  g469(.A1(new_n656), .A2(new_n519), .A3(new_n438), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT46), .Z(new_n672));
  OAI21_X1  g471(.A(G36gat), .B1(new_n668), .B2(new_n375), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(G1329gat));
  INV_X1    g473(.A(G43gat), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n652), .A2(new_n675), .A3(new_n428), .A4(new_n655), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n677), .A2(new_n678), .B1(KEYINPUT104), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n681));
  OAI21_X1  g480(.A(G43gat), .B1(new_n668), .B2(new_n429), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(G1330gat));
  AND2_X1   g484(.A1(new_n656), .A2(new_n471), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G50gat), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n667), .A2(G50gat), .A3(new_n471), .A4(new_n655), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT48), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1331gat));
  AND3_X1   g492(.A1(new_n474), .A2(new_n661), .A3(new_n660), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n662), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n626), .A2(new_n586), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(new_n566), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n310), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT105), .B(G57gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1332gat));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n375), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  AND2_X1   g502(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n702), .B2(new_n703), .ZN(G1333gat));
  INV_X1    g505(.A(G71gat), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n698), .A2(new_n707), .A3(new_n429), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT106), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n428), .B(KEYINPUT107), .Z(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n698), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT50), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n709), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1334gat));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n256), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g517(.A1(new_n696), .A2(new_n514), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n667), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n310), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n474), .A2(new_n661), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n514), .A2(new_n654), .A3(new_n565), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n725), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n626), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n532), .A3(new_n629), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n722), .A2(new_n731), .ZN(G1336gat));
  INV_X1    g531(.A(G92gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n733), .A3(new_n438), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(KEYINPUT52), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n719), .B1(new_n659), .B2(new_n666), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n438), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n531), .A2(new_n533), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n738), .A2(new_n739), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n736), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n738), .A2(new_n741), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT52), .B1(new_n745), .B2(new_n735), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n721), .B2(new_n429), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n535), .A3(new_n428), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT109), .Z(G1338gat));
  AOI21_X1  g550(.A(new_n536), .B1(new_n737), .B2(new_n471), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n256), .A2(G106gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n730), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT51), .B1(new_n723), .B2(new_n725), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n727), .B(new_n724), .C1(new_n474), .C2(new_n661), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n653), .B(new_n754), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT53), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n664), .B1(new_n475), .B2(new_n565), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n565), .A2(new_n664), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n694), .A2(new_n662), .A3(new_n765), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n471), .B(new_n720), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  AOI211_X1 g566(.A(KEYINPUT111), .B(new_n763), .C1(G106gat), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(new_n763), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n761), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n761), .B(KEYINPUT112), .C1(new_n768), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1339gat));
  NAND3_X1  g576(.A1(new_n566), .A2(new_n654), .A3(new_n626), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n603), .A2(new_n589), .A3(new_n604), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n614), .A2(KEYINPUT54), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n782), .B(new_n611), .C1(new_n605), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n613), .A2(new_n783), .A3(new_n588), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT113), .B1(new_n785), .B2(new_n617), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT55), .B(new_n781), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n623), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT54), .B(new_n589), .C1(new_n603), .C2(new_n604), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n789), .B2(new_n611), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(KEYINPUT113), .A3(new_n617), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT55), .B1(new_n792), .B2(new_n781), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n779), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n781), .B1(new_n784), .B2(new_n786), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n623), .A4(new_n787), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n586), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n574), .A2(new_n575), .A3(new_n578), .A4(new_n585), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n576), .A2(new_n577), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n569), .B1(new_n567), .B2(new_n571), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n584), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n800), .B(new_n803), .C1(new_n624), .C2(new_n625), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n565), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n803), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n562), .B2(new_n564), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n794), .A2(new_n807), .A3(new_n798), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT115), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n514), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n805), .A2(KEYINPUT115), .A3(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n778), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n310), .A2(new_n438), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n472), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(new_n257), .A3(new_n654), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n629), .A3(new_n467), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n804), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n651), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n808), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n514), .A3(new_n810), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n310), .B1(new_n823), .B2(new_n778), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(new_n467), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n438), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n586), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n816), .B1(new_n828), .B2(new_n257), .ZN(G1340gat));
  OAI21_X1  g628(.A(G120gat), .B1(new_n815), .B2(new_n626), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT117), .Z(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n258), .A3(new_n653), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n824), .A2(new_n825), .A3(new_n467), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n825), .B1(new_n824), .B2(new_n467), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n375), .B(new_n513), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n827), .B2(new_n513), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n834), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  OAI21_X1  g641(.A(G127gat), .B1(new_n815), .B2(new_n514), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n818), .A2(new_n826), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n839), .A3(new_n375), .A4(new_n513), .ZN(new_n847));
  AOI21_X1  g646(.A(G127gat), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n843), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT119), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n850), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n438), .A2(new_n651), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n846), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n815), .B2(new_n651), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n814), .A2(new_n429), .ZN(new_n859));
  INV_X1    g658(.A(new_n795), .ZN(new_n860));
  XNOR2_X1  g659(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n586), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n804), .B1(new_n788), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n651), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n513), .B1(new_n864), .B2(new_n808), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(KEYINPUT121), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n778), .B1(new_n865), .B2(KEYINPUT121), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n471), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n859), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n256), .B1(new_n823), .B2(new_n778), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n654), .ZN(new_n874));
  INV_X1    g673(.A(new_n859), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n876), .A2(G141gat), .A3(new_n654), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT58), .ZN(G1344gat));
  NOR3_X1   g678(.A1(new_n876), .A2(G148gat), .A3(new_n626), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n869), .A2(new_n872), .A3(new_n653), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(G148gat), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n813), .A2(new_n471), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n788), .A2(new_n793), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n863), .A2(new_n651), .B1(new_n887), .B2(new_n807), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n778), .B1(new_n888), .B2(new_n513), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n256), .A2(KEYINPUT57), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n886), .A2(KEYINPUT57), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n653), .A3(new_n875), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n883), .B1(new_n892), .B2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n881), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n896), .B(new_n881), .C1(new_n885), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1345gat));
  OAI21_X1  g697(.A(G155gat), .B1(new_n873), .B2(new_n514), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n513), .A2(new_n206), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n876), .B2(new_n900), .ZN(G1346gat));
  OAI21_X1  g700(.A(G162gat), .B1(new_n873), .B2(new_n651), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n256), .A2(G162gat), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n824), .A2(new_n429), .A3(new_n853), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n905), .B(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n629), .A2(new_n375), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n813), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(new_n467), .ZN(new_n910));
  AOI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n586), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n710), .A2(new_n471), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(G169gat), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n654), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n911), .A2(new_n915), .ZN(G1348gat));
  INV_X1    g715(.A(G176gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n910), .A2(new_n917), .A3(new_n653), .ZN(new_n918));
  OAI21_X1  g717(.A(G176gat), .B1(new_n913), .B2(new_n626), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT124), .Z(G1349gat));
  OAI211_X1 g720(.A(new_n910), .B(new_n513), .C1(new_n347), .C2(new_n346), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n325), .B1(new_n913), .B2(new_n514), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n922), .A2(new_n923), .B1(KEYINPUT125), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT125), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n913), .B2(new_n651), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT61), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n333), .A3(new_n565), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1351gat));
  NAND2_X1  g730(.A1(new_n908), .A2(new_n429), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n886), .A2(G197gat), .A3(new_n654), .A4(new_n932), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT126), .Z(new_n934));
  NAND2_X1  g733(.A1(new_n889), .A2(new_n890), .ZN(new_n935));
  INV_X1    g734(.A(new_n932), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n936), .C1(new_n870), .C2(new_n871), .ZN(new_n937));
  OAI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n654), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(G1352gat));
  NOR4_X1   g738(.A1(new_n886), .A2(G204gat), .A3(new_n626), .A4(new_n932), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n891), .A2(new_n653), .A3(new_n936), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G204gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1353gat));
  NOR2_X1   g743(.A1(new_n886), .A2(new_n932), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n227), .A3(new_n513), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n937), .A2(new_n514), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n227), .B1(new_n947), .B2(KEYINPUT127), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(KEYINPUT63), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n937), .B2(new_n651), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n945), .A2(new_n228), .A3(new_n565), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1355gat));
endmodule


