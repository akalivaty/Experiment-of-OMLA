

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U323 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U324 ( .A(n555), .B(KEYINPUT74), .ZN(n560) );
  XOR2_X1 U325 ( .A(n318), .B(n317), .Z(n290) );
  XNOR2_X1 U326 ( .A(n386), .B(n385), .ZN(n529) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT114), .ZN(n403) );
  XNOR2_X1 U328 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U329 ( .A(KEYINPUT87), .ZN(n445) );
  XNOR2_X1 U330 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n385) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U332 ( .A(n319), .B(n290), .ZN(n320) );
  XNOR2_X1 U333 ( .A(n367), .B(n366), .ZN(n368) );
  INV_X1 U334 ( .A(KEYINPUT100), .ZN(n471) );
  XNOR2_X1 U335 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U336 ( .A(n369), .B(n368), .ZN(n379) );
  XNOR2_X1 U337 ( .A(n471), .B(KEYINPUT38), .ZN(n472) );
  XNOR2_X1 U338 ( .A(n473), .B(n472), .ZN(n500) );
  XNOR2_X1 U339 ( .A(G183GAT), .B(KEYINPUT120), .ZN(n455) );
  XNOR2_X1 U340 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n474) );
  XNOR2_X1 U341 ( .A(n456), .B(n455), .ZN(G1350GAT) );
  XNOR2_X1 U342 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n292) );
  XNOR2_X1 U344 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n308) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n358) );
  XOR2_X1 U347 ( .A(G134GAT), .B(G99GAT), .Z(n294) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(n358), .B(n295), .Z(n297) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G15GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U356 ( .A(n301), .B(n300), .Z(n306) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n302), .B(G127GAT), .ZN(n407) );
  XOR2_X1 U359 ( .A(G183GAT), .B(KEYINPUT19), .Z(n304) );
  XNOR2_X1 U360 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n398) );
  XNOR2_X1 U362 ( .A(n407), .B(n398), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U364 ( .A(n308), .B(n307), .Z(n522) );
  INV_X1 U365 ( .A(n522), .ZN(n530) );
  INV_X1 U366 ( .A(KEYINPUT47), .ZN(n376) );
  XOR2_X1 U367 ( .A(KEYINPUT7), .B(G50GAT), .Z(n310) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G29GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U370 ( .A(KEYINPUT8), .B(n311), .Z(n349) );
  XOR2_X1 U371 ( .A(G92GAT), .B(KEYINPUT73), .Z(n313) );
  XNOR2_X1 U372 ( .A(G190GAT), .B(G218GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U374 ( .A(G36GAT), .B(n314), .Z(n393) );
  XNOR2_X1 U375 ( .A(n349), .B(n393), .ZN(n323) );
  XOR2_X1 U376 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n316) );
  XOR2_X1 U377 ( .A(G134GAT), .B(KEYINPUT72), .Z(n419) );
  XOR2_X1 U378 ( .A(G99GAT), .B(G85GAT), .Z(n363) );
  XNOR2_X1 U379 ( .A(n419), .B(n363), .ZN(n315) );
  XNOR2_X1 U380 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U381 ( .A(G162GAT), .B(G106GAT), .Z(n437) );
  XNOR2_X1 U382 ( .A(n437), .B(KEYINPUT71), .ZN(n319) );
  XOR2_X1 U383 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n318) );
  NAND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n555) );
  XOR2_X1 U386 ( .A(G78GAT), .B(G211GAT), .Z(n325) );
  XNOR2_X1 U387 ( .A(G127GAT), .B(G71GAT), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U389 ( .A(n326), .B(G155GAT), .Z(n328) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G1GAT), .Z(n342) );
  XNOR2_X1 U391 ( .A(n342), .B(G22GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n333) );
  XNOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n329), .B(KEYINPUT13), .ZN(n361) );
  XOR2_X1 U395 ( .A(n361), .B(G64GAT), .Z(n331) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U399 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n335) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(KEYINPUT15), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U402 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n337) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U406 ( .A(n341), .B(n340), .Z(n575) );
  INV_X1 U407 ( .A(n575), .ZN(n537) );
  XOR2_X1 U408 ( .A(G169GAT), .B(G8GAT), .Z(n399) );
  XNOR2_X1 U409 ( .A(n342), .B(n399), .ZN(n353) );
  XOR2_X1 U410 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n344) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U413 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XOR2_X1 U414 ( .A(n345), .B(n439), .Z(n351) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(G113GAT), .Z(n347) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G197GAT), .ZN(n346) );
  XNOR2_X1 U417 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n568) );
  XNOR2_X1 U421 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n355) );
  AND2_X1 U422 ( .A1(G230GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n357) );
  INV_X1 U424 ( .A(KEYINPUT33), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n360) );
  XOR2_X1 U426 ( .A(G176GAT), .B(G64GAT), .Z(n396) );
  XNOR2_X1 U427 ( .A(n358), .B(n396), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U429 ( .A(n362), .B(n361), .Z(n369) );
  XOR2_X1 U430 ( .A(G148GAT), .B(G78GAT), .Z(n436) );
  XNOR2_X1 U431 ( .A(n436), .B(n363), .ZN(n367) );
  XOR2_X1 U432 ( .A(KEYINPUT69), .B(G92GAT), .Z(n365) );
  XNOR2_X1 U433 ( .A(G204GAT), .B(G106GAT), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U435 ( .A(KEYINPUT41), .B(n379), .Z(n550) );
  NOR2_X1 U436 ( .A1(n568), .A2(n550), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n370), .B(KEYINPUT46), .ZN(n371) );
  NOR2_X1 U438 ( .A1(n537), .A2(n371), .ZN(n373) );
  INV_X1 U439 ( .A(KEYINPUT108), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U441 ( .A1(n555), .A2(n374), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n568), .B(KEYINPUT67), .ZN(n558) );
  XNOR2_X1 U444 ( .A(KEYINPUT36), .B(n560), .ZN(n580) );
  NAND2_X1 U445 ( .A1(n537), .A2(n580), .ZN(n378) );
  XNOR2_X1 U446 ( .A(KEYINPUT45), .B(KEYINPUT109), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n378), .B(n377), .ZN(n380) );
  NAND2_X1 U448 ( .A1(n380), .A2(n379), .ZN(n381) );
  NOR2_X1 U449 ( .A1(n558), .A2(n381), .ZN(n382) );
  XNOR2_X1 U450 ( .A(KEYINPUT110), .B(n382), .ZN(n383) );
  NOR2_X1 U451 ( .A1(n384), .A2(n383), .ZN(n386) );
  XOR2_X1 U452 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n388) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U455 ( .A(n389), .B(KEYINPUT93), .Z(n395) );
  XOR2_X1 U456 ( .A(KEYINPUT84), .B(G211GAT), .Z(n391) );
  XNOR2_X1 U457 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U459 ( .A(G197GAT), .B(n392), .Z(n449) );
  XNOR2_X1 U460 ( .A(n449), .B(n393), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U462 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U464 ( .A(n401), .B(n400), .Z(n507) );
  XNOR2_X1 U465 ( .A(KEYINPUT113), .B(n507), .ZN(n402) );
  NOR2_X1 U466 ( .A1(n529), .A2(n402), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n428) );
  XOR2_X1 U468 ( .A(G155GAT), .B(KEYINPUT85), .Z(n406) );
  XNOR2_X1 U469 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n444) );
  XNOR2_X1 U471 ( .A(n407), .B(n444), .ZN(n427) );
  XOR2_X1 U472 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n409) );
  XNOR2_X1 U473 ( .A(G120GAT), .B(G148GAT), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U475 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n411) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G57GAT), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U478 ( .A(n413), .B(n412), .Z(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n415) );
  XNOR2_X1 U480 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n423) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G162GAT), .Z(n417) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G141GAT), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U485 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U490 ( .A(n427), .B(n426), .Z(n545) );
  INV_X1 U491 ( .A(n545), .ZN(n518) );
  NAND2_X1 U492 ( .A1(n428), .A2(n518), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n429), .B(KEYINPUT65), .ZN(n565) );
  XOR2_X1 U494 ( .A(KEYINPUT82), .B(KEYINPUT86), .Z(n431) );
  XNOR2_X1 U495 ( .A(G50GAT), .B(G218GAT), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT83), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U498 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U500 ( .A(n435), .B(n434), .Z(n443) );
  XOR2_X1 U501 ( .A(n437), .B(n436), .Z(n441) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n444), .B(KEYINPUT88), .ZN(n446) );
  XOR2_X1 U505 ( .A(n450), .B(n449), .Z(n462) );
  NAND2_X1 U506 ( .A1(n565), .A2(n462), .ZN(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT55), .B(KEYINPUT115), .Z(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U509 ( .A1(n530), .A2(n453), .ZN(n454) );
  XOR2_X2 U510 ( .A(KEYINPUT116), .B(n454), .Z(n561) );
  NAND2_X1 U511 ( .A1(n561), .A2(n537), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n507), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U513 ( .A1(n530), .A2(n462), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U515 ( .A1(n463), .A2(n566), .ZN(n544) );
  NAND2_X1 U516 ( .A1(n530), .A2(n507), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n462), .A2(n458), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n459), .Z(n460) );
  NAND2_X1 U519 ( .A1(n544), .A2(n460), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n461), .A2(n518), .ZN(n467) );
  XOR2_X1 U521 ( .A(n462), .B(KEYINPUT28), .Z(n513) );
  INV_X1 U522 ( .A(n513), .ZN(n525) );
  NAND2_X1 U523 ( .A1(n463), .A2(n525), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n518), .A2(n464), .ZN(n531) );
  XNOR2_X1 U525 ( .A(n531), .B(KEYINPUT96), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n465), .A2(n522), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n483) );
  NAND2_X1 U528 ( .A1(n575), .A2(n483), .ZN(n468) );
  XNOR2_X1 U529 ( .A(KEYINPUT99), .B(n468), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n469), .A2(n580), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT37), .B(n470), .Z(n517) );
  NAND2_X1 U532 ( .A1(n558), .A2(n379), .ZN(n485) );
  NOR2_X1 U533 ( .A1(n517), .A2(n485), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n518), .A2(n500), .ZN(n475) );
  INV_X1 U535 ( .A(n550), .ZN(n534) );
  NAND2_X1 U536 ( .A1(n534), .A2(n561), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n477) );
  XNOR2_X1 U538 ( .A(KEYINPUT117), .B(KEYINPUT57), .ZN(n476) );
  XOR2_X1 U539 ( .A(n477), .B(n476), .Z(n479) );
  XOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT56), .Z(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1349GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n487) );
  NOR2_X1 U544 ( .A1(n575), .A2(n560), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n482), .B(KEYINPUT16), .ZN(n484) );
  NAND2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n503) );
  NOR2_X1 U547 ( .A1(n485), .A2(n503), .ZN(n493) );
  NAND2_X1 U548 ( .A1(n493), .A2(n545), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n507), .A2(n493), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n491) );
  NAND2_X1 U554 ( .A1(n493), .A2(n530), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n493), .A2(n513), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 U559 ( .A(n507), .ZN(n520) );
  NOR2_X1 U560 ( .A1(n520), .A2(n500), .ZN(n495) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n497) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n497), .B(n496), .ZN(n499) );
  NOR2_X1 U565 ( .A1(n522), .A2(n500), .ZN(n498) );
  XOR2_X1 U566 ( .A(n499), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U567 ( .A1(n525), .A2(n500), .ZN(n501) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NAND2_X1 U569 ( .A1(n534), .A2(n568), .ZN(n502) );
  XOR2_X1 U570 ( .A(KEYINPUT103), .B(n502), .Z(n516) );
  NOR2_X1 U571 ( .A1(n516), .A2(n503), .ZN(n504) );
  XNOR2_X1 U572 ( .A(KEYINPUT104), .B(n504), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n512), .A2(n545), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n509) );
  NAND2_X1 U577 ( .A1(n512), .A2(n507), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n512), .A2(n530), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  OR2_X1 U585 ( .A1(n517), .A2(n516), .ZN(n524) );
  NOR2_X1 U586 ( .A1(n518), .A2(n524), .ZN(n519) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n520), .A2(n524), .ZN(n521) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n522), .A2(n524), .ZN(n523) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT107), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n529), .A2(n532), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n558), .A2(n540), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U601 ( .A1(n540), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n540), .A2(n537), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT51), .B(KEYINPUT111), .Z(n542) );
  NAND2_X1 U607 ( .A1(n540), .A2(n560), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NOR2_X1 U610 ( .A1(n529), .A2(n544), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n568), .A2(n554), .ZN(n547) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT112), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n550), .A2(n554), .ZN(n551) );
  XOR2_X1 U618 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NOR2_X1 U619 ( .A1(n575), .A2(n554), .ZN(n553) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  INV_X1 U621 ( .A(n554), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U631 ( .A(n567), .B(KEYINPUT122), .Z(n581) );
  INV_X1 U632 ( .A(n581), .ZN(n576) );
  NOR2_X1 U633 ( .A1(n576), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n576), .A2(n379), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT124), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1355GAT) );
endmodule

