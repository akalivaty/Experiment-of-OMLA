//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n438, new_n439, new_n440, new_n443, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n438));
  OR2_X1    g013(.A1(new_n438), .A2(G69), .ZN(new_n439));
  NAND2_X1  g014(.A1(new_n438), .A2(G69), .ZN(new_n440));
  NAND2_X1  g015(.A1(new_n439), .A2(new_n440), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G57), .Z(new_n443));
  INV_X1    g018(.A(new_n443), .ZN(G237));
  INV_X1    g019(.A(G108), .ZN(G238));
  NAND4_X1  g020(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT70), .ZN(G319));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n469), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n473));
  OR2_X1    g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NOR2_X1   g064(.A1(new_n477), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G102), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n469), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n471), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n478), .A2(new_n480), .A3(G138), .A4(new_n471), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n471), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n503), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n510), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n505), .A2(new_n506), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n514), .A2(G51), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n523), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n522), .A2(G90), .B1(G52), .B2(new_n514), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n521), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n509), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n514), .A2(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n517), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(new_n514), .A2(G53), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT9), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n522), .A2(G91), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n550), .B(new_n551), .C1(new_n509), .C2(new_n552), .ZN(G299));
  NAND2_X1  g128(.A1(G171), .A2(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n530), .A2(new_n534), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  NAND3_X1  g135(.A1(new_n507), .A2(G87), .A3(new_n516), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n522), .A2(new_n563), .A3(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n514), .A2(G49), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  AND3_X1   g143(.A1(new_n505), .A2(G61), .A3(new_n506), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n505), .A2(G86), .A3(new_n506), .ZN(new_n573));
  NAND2_X1  g148(.A1(G48), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(new_n516), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n522), .A2(G85), .B1(G47), .B2(new_n514), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n509), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(new_n522), .A2(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n514), .A2(G54), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n509), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n558), .B2(new_n591), .ZN(G284));
  OAI21_X1  g168(.A(new_n592), .B1(new_n558), .B2(new_n591), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  AND3_X1   g173(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n599));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n482), .A2(G123), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT77), .Z(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n609), .B(new_n610), .C1(G111), .C2(new_n471), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n484), .A2(G135), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2096), .Z(new_n614));
  NAND2_X1  g189(.A1(new_n469), .A2(new_n490), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(KEYINPUT76), .B2(G2100), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT76), .B(G2100), .Z(new_n619));
  OAI211_X1 g194(.A(new_n614), .B(new_n618), .C1(new_n617), .C2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2443), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n631), .B(new_n632), .Z(new_n633));
  AND2_X1   g208(.A1(new_n633), .A2(G14), .ZN(G401));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2072), .B(G2078), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT18), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(KEYINPUT17), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n643), .A2(new_n636), .A3(new_n639), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n639), .B1(new_n637), .B2(new_n642), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n638), .B(KEYINPUT81), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n637), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n652), .A2(new_n653), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n658), .A2(new_n654), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n663), .ZN(new_n666));
  NAND4_X1  g241(.A1(new_n662), .A2(new_n664), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G24), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n580), .A2(new_n582), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n675), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(KEYINPUT91), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(G23), .ZN(new_n683));
  INV_X1    g258(.A(G288), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n675), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT33), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT89), .B1(new_n689), .B2(G16), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n689), .A2(KEYINPUT89), .A3(G16), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(G166), .C2(new_n675), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT90), .B(G1971), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n675), .A2(G6), .ZN(new_n695));
  INV_X1    g270(.A(G305), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n675), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n688), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n682), .B1(KEYINPUT34), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n482), .A2(G119), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n484), .A2(G131), .ZN(new_n703));
  NOR2_X1   g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(KEYINPUT85), .A2(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(KEYINPUT85), .A2(G29), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(new_n706), .B(G25), .S(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  OR2_X1    g289(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n701), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n716), .A2(KEYINPUT91), .A3(new_n681), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G139), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n718), .B(new_n721), .C1(new_n471), .C2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  MUX2_X1   g299(.A(G33), .B(new_n724), .S(G29), .Z(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G2072), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT98), .B(KEYINPUT31), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G11), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT24), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(G34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(G34), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n709), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n475), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  NOR2_X1   g312(.A1(G164), .A2(new_n709), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G27), .B2(new_n709), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT30), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n613), .B2(new_n709), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n733), .A2(G32), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n482), .A2(G129), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n484), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n490), .A2(G105), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND4_X1  g325(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n745), .B1(new_n752), .B2(new_n733), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n756), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n744), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n726), .A2(new_n728), .A3(new_n740), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n739), .A2(new_n737), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n675), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n675), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1961), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G21), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G168), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1966), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n725), .A2(G2072), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT96), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n765), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT99), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n681), .A2(KEYINPUT91), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n701), .A2(new_n774), .A3(new_n714), .A4(new_n715), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n542), .B2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1341), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n675), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n599), .B2(new_n675), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n709), .A2(G35), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G162), .B2(new_n709), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT29), .ZN(new_n785));
  INV_X1    g360(.A(G2090), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n675), .A2(G20), .ZN(new_n788));
  OAI211_X1 g363(.A(KEYINPUT23), .B(new_n788), .C1(new_n596), .C2(new_n675), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(KEYINPUT23), .B2(new_n788), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n778), .A2(new_n782), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n772), .B2(KEYINPUT99), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n717), .A2(new_n773), .A3(new_n775), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n484), .A2(G140), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n482), .A2(G128), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n471), .A2(G116), .ZN(new_n797));
  OR3_X1    g372(.A1(KEYINPUT92), .A2(G104), .A3(G2105), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT92), .B1(G104), .B2(G2105), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n798), .A2(G2104), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n709), .A2(G26), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT94), .B(G2067), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n794), .A2(new_n808), .ZN(G311));
  INV_X1    g384(.A(G311), .ZN(G150));
  XOR2_X1   g385(.A(KEYINPUT101), .B(G55), .Z(new_n811));
  AOI22_X1  g386(.A1(new_n522), .A2(G93), .B1(new_n514), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n509), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT102), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n600), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT39), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n542), .A2(new_n814), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n541), .A2(new_n814), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n819), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n817), .B1(new_n826), .B2(G860), .ZN(G145));
  XNOR2_X1  g402(.A(new_n801), .B(new_n751), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n498), .A2(KEYINPUT103), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n496), .A2(new_n497), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n493), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n828), .B(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(new_n723), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n484), .A2(G142), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n482), .A2(G130), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n839), .B1(new_n836), .B2(new_n835), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n706), .B(new_n616), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n833), .A2(new_n724), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n834), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n834), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(KEYINPUT105), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n834), .A2(new_n849), .A3(new_n844), .A4(new_n845), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n613), .B(G160), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n488), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  INV_X1    g429(.A(new_n846), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n847), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n853), .B(new_n854), .C1(new_n856), .C2(new_n852), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g433(.A1(new_n814), .A2(new_n591), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n677), .A2(G303), .ZN(new_n860));
  NAND2_X1  g435(.A1(G290), .A2(G166), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(G305), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(G305), .B1(new_n860), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(G288), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n684), .A3(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT42), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n821), .B1(new_n542), .B2(new_n814), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n602), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n599), .A2(new_n596), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n590), .A2(G299), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT41), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n874), .B2(new_n871), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n869), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n859), .B1(new_n878), .B2(new_n591), .ZN(G295));
  OAI21_X1  g454(.A(new_n859), .B1(new_n878), .B2(new_n591), .ZN(G331));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n558), .B2(G286), .ZN(new_n882));
  AOI21_X1  g457(.A(G286), .B1(new_n554), .B2(new_n557), .ZN(new_n883));
  NOR2_X1   g458(.A1(G168), .A2(new_n555), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT106), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n823), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n870), .A2(new_n885), .A3(new_n882), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(KEYINPUT107), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n890), .A3(new_n823), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n874), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n874), .B(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n887), .B2(new_n888), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n896), .B2(new_n868), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n865), .A2(new_n867), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n892), .B2(new_n895), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT43), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n892), .A2(new_n898), .A3(new_n895), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n889), .A2(new_n875), .A3(new_n891), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n887), .A2(new_n873), .A3(new_n872), .A4(new_n888), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n905));
  NOR4_X1   g480(.A1(new_n901), .A2(new_n904), .A3(new_n905), .A4(G37), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n897), .B2(new_n899), .ZN(new_n909));
  NOR4_X1   g484(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT43), .A4(G37), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(G397));
  NAND2_X1  g487(.A1(G114), .A2(G2104), .ZN(new_n913));
  INV_X1    g488(.A(G126), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n481), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n915), .A2(G2105), .B1(G102), .B2(new_n490), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n496), .A2(new_n497), .A3(new_n830), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n830), .B1(new_n496), .B2(new_n497), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT45), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n472), .A2(new_n474), .A3(G40), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(G1996), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT108), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(new_n751), .ZN(new_n926));
  INV_X1    g501(.A(G2067), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n801), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT109), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n929), .B2(new_n752), .ZN(new_n930));
  INV_X1    g505(.A(G1996), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OR3_X1    g508(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT110), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT110), .B1(new_n926), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n706), .A2(new_n713), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n706), .A2(new_n713), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n921), .B(new_n922), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n677), .A2(new_n679), .ZN(new_n941));
  NAND2_X1  g516(.A1(G290), .A2(G1986), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n923), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n936), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n919), .A2(KEYINPUT45), .A3(new_n920), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n920), .B1(new_n493), .B2(new_n498), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n945), .A2(new_n737), .A3(new_n922), .A4(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  INV_X1    g527(.A(G1961), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n832), .B2(G1384), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n919), .A2(KEYINPUT111), .A3(new_n920), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT50), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n946), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n922), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT124), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n949), .A2(new_n962), .A3(new_n950), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n945), .A2(new_n922), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n950), .A2(G2078), .ZN(new_n965));
  INV_X1    g540(.A(new_n921), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n952), .A2(new_n961), .A3(new_n963), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G171), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n949), .A2(new_n962), .A3(new_n950), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n962), .B1(new_n949), .B2(new_n950), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n955), .A2(new_n947), .A3(new_n956), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n922), .A3(new_n965), .A4(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n972), .A2(G301), .A3(new_n975), .A4(new_n961), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n969), .A2(new_n976), .A3(KEYINPUT54), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n922), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n768), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n955), .A2(new_n956), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n959), .ZN(new_n981));
  INV_X1    g556(.A(new_n960), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n735), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT112), .B(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(G286), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n979), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n960), .B1(new_n980), .B2(new_n959), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n768), .A2(new_n978), .B1(new_n987), .B2(new_n735), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(G8), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n986), .B(KEYINPUT51), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n992));
  INV_X1    g567(.A(new_n984), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n992), .B(new_n985), .C1(new_n988), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n996));
  NAND4_X1  g571(.A1(new_n952), .A2(new_n961), .A3(new_n963), .A4(new_n975), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n558), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n972), .A2(G301), .A3(new_n961), .A4(new_n967), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n977), .A2(new_n995), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n572), .B2(new_n576), .ZN(new_n1005));
  OR3_X1    g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n832), .A2(new_n954), .A3(G1384), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT111), .B1(new_n919), .B2(new_n920), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n922), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n1009), .A3(new_n984), .A4(new_n1010), .ZN(new_n1011));
  AND4_X1   g586(.A1(G1976), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1013), .A2(new_n1009), .A3(new_n984), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n922), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n955), .B2(new_n956), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1018), .A2(new_n993), .A3(new_n1012), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1011), .B(new_n1016), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT114), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1009), .A2(new_n984), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n1023), .B2(new_n1012), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1011), .A4(new_n1016), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n945), .A2(new_n922), .A3(new_n948), .ZN(new_n1028));
  INV_X1    g603(.A(G1971), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n958), .A2(new_n959), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n922), .B(new_n1031), .C1(new_n980), .C2(new_n959), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1032), .B2(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n984), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n510), .B2(new_n519), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT55), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n981), .A2(new_n786), .A3(new_n982), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1030), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1036), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  AND4_X1   g616(.A1(KEYINPUT125), .A2(new_n1027), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n1043), .B(new_n1036), .C1(new_n1038), .C2(new_n1030), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT125), .B1(new_n1045), .B2(new_n1037), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1001), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1956), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1032), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n964), .A2(new_n948), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n550), .B2(KEYINPUT115), .ZN(new_n1052));
  XNOR2_X1  g627(.A(G299), .B(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT58), .B(G1341), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT119), .B(G1996), .Z(new_n1059));
  OAI22_X1  g634(.A1(new_n1018), .A2(new_n1058), .B1(new_n1028), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n542), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(KEYINPUT59), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(KEYINPUT59), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT120), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1057), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT116), .B1(new_n1009), .B2(G2067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n781), .B1(new_n957), .B2(new_n960), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1018), .A2(new_n1070), .A3(new_n927), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1068), .A2(new_n1069), .A3(new_n1074), .A4(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n590), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1056), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT122), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(new_n1056), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(KEYINPUT60), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(new_n1084), .A3(new_n1075), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n599), .A3(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1067), .A2(new_n1077), .A3(new_n1082), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1073), .A2(new_n599), .A3(new_n1075), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1055), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1054), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1047), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1011), .A2(new_n1014), .A3(new_n684), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1002), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g671(.A(KEYINPUT113), .B1(new_n1041), .B2(new_n1021), .C1(new_n1096), .C2(new_n1023), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1041), .A2(new_n1021), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1023), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n988), .A2(G286), .A3(new_n993), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1043), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1040), .B2(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1044), .A2(new_n1021), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT63), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1045), .A2(new_n1108), .A3(new_n1037), .A4(new_n1103), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1102), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n991), .A2(new_n994), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n998), .B1(new_n1111), .B2(KEYINPUT62), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n995), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(new_n1114), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n944), .B1(new_n1093), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n801), .A2(G2067), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n923), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n941), .A2(new_n923), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT48), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n936), .A2(new_n940), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT46), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n925), .B(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n930), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1120), .A2(new_n1123), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1117), .A2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g708(.A1(G401), .A2(G227), .ZN(new_n1135));
  NAND2_X1  g709(.A1(new_n1135), .A2(new_n857), .ZN(new_n1136));
  INV_X1    g710(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g711(.A(G319), .ZN(new_n1138));
  OR2_X1    g712(.A1(new_n1138), .A2(G229), .ZN(new_n1139));
  INV_X1    g713(.A(new_n1139), .ZN(new_n1140));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1140), .C1(new_n909), .C2(new_n910), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


