//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G128), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n200), .A2(G137), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n200), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .A4(new_n201), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n194), .B(new_n196), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n199), .A2(new_n204), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n206), .A2(new_n208), .A3(new_n201), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n215), .A2(new_n210), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT0), .B(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT64), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n194), .A2(new_n196), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n197), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n219), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n213), .B1(new_n216), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT2), .B(G113), .Z(new_n229));
  XNOR2_X1  g043(.A(G116), .B(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(new_n230), .B(KEYINPUT66), .Z(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n229), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT30), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(KEYINPUT65), .A3(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT30), .B(new_n213), .C1(new_n216), .C2(new_n227), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n241), .A2(new_n233), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n217), .A2(new_n218), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n221), .B1(new_n244), .B2(new_n225), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n215), .A2(new_n210), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n219), .ZN(new_n247));
  AOI211_X1 g061(.A(new_n237), .B(KEYINPUT30), .C1(new_n247), .C2(new_n213), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT65), .B1(new_n228), .B2(new_n235), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n242), .B(KEYINPUT67), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n192), .B(new_n234), .C1(new_n243), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n228), .A2(new_n233), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n228), .A2(new_n233), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(KEYINPUT28), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n255), .A2(KEYINPUT28), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n192), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT29), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n234), .A2(new_n261), .A3(new_n253), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n228), .A2(new_n233), .A3(KEYINPUT68), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT28), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n264), .A2(KEYINPUT29), .A3(new_n191), .A4(new_n257), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(G472), .B1(new_n260), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n270), .B(G472), .C1(new_n260), .C2(new_n267), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n255), .A2(new_n192), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n243), .B2(new_n251), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n256), .A2(new_n257), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n192), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n242), .B1(new_n248), .B2(new_n249), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n250), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT31), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n272), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NOR2_X1   g098(.A1(G472), .A2(G902), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n269), .B(new_n271), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT9), .B(G234), .ZN(new_n289));
  OAI21_X1  g103(.A(G221), .B1(new_n289), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n293));
  INV_X1    g107(.A(G104), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(G107), .ZN(new_n295));
  INV_X1    g109(.A(G107), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT3), .A3(G104), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G101), .ZN(new_n299));
  OR3_X1    g113(.A1(new_n296), .A2(KEYINPUT73), .A3(G104), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(G107), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n294), .B2(G107), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n296), .A3(G104), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n306), .A3(new_n301), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G101), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n303), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n292), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n303), .A2(new_n308), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT76), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(KEYINPUT77), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n199), .A2(new_n212), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT10), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n298), .A2(new_n302), .A3(new_n300), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G101), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n303), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n227), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n322), .B(G101), .C1(new_n324), .C2(new_n325), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n319), .B1(new_n313), .B2(new_n318), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n216), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n320), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n312), .B2(new_n316), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n246), .B1(new_n336), .B2(new_n332), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G140), .ZN(new_n338));
  INV_X1    g152(.A(G227), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G953), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n334), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OR2_X1    g158(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n345));
  INV_X1    g159(.A(new_n318), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n310), .A2(new_n311), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n313), .A2(new_n318), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n246), .B(new_n345), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n314), .A2(new_n318), .A3(new_n315), .ZN(new_n350));
  INV_X1    g164(.A(new_n348), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n216), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n353));
  OAI21_X1  g167(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n342), .B1(new_n334), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT79), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n334), .A2(new_n354), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n357), .B(new_n343), .C1(new_n358), .C2(new_n342), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n359), .A3(G469), .ZN(new_n360));
  INV_X1    g174(.A(G469), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n266), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n216), .B1(new_n321), .B2(new_n333), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n336), .A2(new_n246), .A3(new_n332), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n341), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n334), .A2(new_n354), .A3(new_n342), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n362), .B1(new_n367), .B2(new_n361), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n291), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G953), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n370), .A2(G952), .ZN(new_n371));
  NAND2_X1  g185(.A1(G234), .A2(G237), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(G902), .A3(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT21), .B(G898), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G214), .B1(G237), .B2(G902), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n379), .B(KEYINPUT80), .Z(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G210), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G125), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n318), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n328), .B2(new_n384), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n370), .A2(G224), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G122), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n389), .B(KEYINPUT81), .Z(new_n390));
  INV_X1    g204(.A(G119), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G116), .ZN(new_n392));
  OAI21_X1  g206(.A(G113), .B1(new_n392), .B2(KEYINPUT5), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n230), .B(KEYINPUT66), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n231), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n312), .B2(new_n316), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n233), .A2(new_n327), .A3(new_n329), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n389), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT6), .B(new_n390), .C1(new_n399), .C2(new_n400), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n388), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n313), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n230), .A2(KEYINPUT5), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(KEYINPUT82), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n393), .B1(new_n409), .B2(KEYINPUT82), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n410), .A2(new_n411), .B1(new_n229), .B2(new_n230), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n413));
  OAI22_X1  g227(.A1(new_n412), .A2(new_n413), .B1(new_n310), .B2(new_n311), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n389), .B(KEYINPUT8), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n387), .A2(KEYINPUT7), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n386), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n266), .B1(new_n423), .B2(new_n403), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n383), .B1(new_n407), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n421), .B1(new_n416), .B2(new_n418), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n397), .A2(new_n231), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n317), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n400), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n389), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n406), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(KEYINPUT6), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n401), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n431), .B(new_n382), .C1(new_n434), .C2(new_n388), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n381), .B1(new_n425), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n369), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n294), .ZN(new_n439));
  XNOR2_X1  g253(.A(G125), .B(G140), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(new_n193), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n442));
  AOI21_X1  g256(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT18), .B(G131), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n187), .A2(G214), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n195), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT18), .A2(G131), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n441), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n384), .A2(KEYINPUT16), .A3(G140), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n440), .B2(KEYINPUT16), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G146), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n193), .B(new_n451), .C1(KEYINPUT16), .C2(new_n440), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  OAI21_X1  g270(.A(G131), .B1(new_n442), .B2(new_n443), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n446), .A2(new_n209), .A3(new_n447), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n457), .A2(new_n459), .A3(new_n456), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n439), .B(new_n450), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G140), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n384), .A2(G140), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT84), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT19), .ZN(new_n468));
  AND4_X1   g282(.A1(new_n463), .A2(new_n464), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT19), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n193), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT85), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n457), .A2(new_n459), .B1(new_n452), .B2(G146), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n193), .C1(new_n469), .C2(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n450), .ZN(new_n478));
  INV_X1    g292(.A(new_n439), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n477), .B1(new_n476), .B2(new_n450), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n461), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n483));
  NOR2_X1   g297(.A1(G475), .A2(G902), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n461), .B(new_n485), .C1(new_n480), .C2(new_n481), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT20), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n491));
  NOR3_X1   g305(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n450), .B1(new_n458), .B2(new_n460), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n495), .A2(new_n479), .ZN(new_n496));
  INV_X1    g310(.A(new_n461), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n266), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G475), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n211), .B2(G143), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n211), .A2(G143), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n195), .A2(G128), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n500), .ZN(new_n505));
  OAI21_X1  g319(.A(G134), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT90), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n502), .A3(new_n200), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT91), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT89), .B1(new_n510), .B2(G116), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n512));
  INV_X1    g326(.A(G116), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(G122), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n513), .A2(G122), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n296), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n296), .B1(new_n515), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n509), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n515), .A2(KEYINPUT14), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n516), .B1(new_n515), .B2(KEYINPUT14), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n296), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n504), .A2(new_n502), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G134), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n508), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n518), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n507), .A2(new_n521), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G217), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n289), .A2(new_n530), .A3(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  OAI221_X1 g347(.A(new_n531), .B1(new_n524), .B2(new_n528), .C1(new_n507), .C2(new_n521), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT92), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G478), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n541), .B2(new_n537), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n494), .A2(new_n499), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n530), .B1(G234), .B2(new_n266), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT22), .B(G137), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n370), .A2(G221), .A3(G234), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n554), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT23), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n391), .B2(G128), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(new_n562), .C1(G119), .C2(new_n211), .ZN(new_n563));
  XNOR2_X1  g377(.A(G119), .B(G128), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  AOI22_X1  g379(.A1(new_n563), .A2(G110), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n453), .B2(new_n454), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT70), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n569), .B(new_n566), .C1(new_n453), .C2(new_n454), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI22_X1  g385(.A1(new_n563), .A2(G110), .B1(new_n564), .B2(new_n565), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n452), .A2(G146), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n440), .A2(new_n193), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n559), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n558), .B(new_n577), .C1(new_n568), .C2(new_n570), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n266), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT25), .B(new_n266), .C1(new_n576), .C2(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n548), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n576), .A2(new_n578), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n584), .A2(G902), .A3(new_n547), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n288), .A2(new_n437), .A3(new_n546), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND2_X1  g402(.A1(new_n283), .A2(new_n285), .ZN(new_n589));
  INV_X1    g403(.A(new_n272), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n279), .B2(new_n250), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT31), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n592), .B2(new_n276), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n589), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n360), .A2(new_n368), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n586), .A3(new_n290), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n379), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n599), .B(new_n377), .C1(new_n425), .C2(new_n435), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n494), .A2(new_n499), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n533), .A2(new_n534), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT33), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n533), .A2(new_n604), .A3(new_n534), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n535), .A2(new_n538), .ZN(new_n608));
  NAND2_X1  g422(.A1(G478), .A2(G902), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n600), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  AND2_X1   g429(.A1(new_n483), .A2(new_n486), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n492), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n490), .A2(new_n491), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n499), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n540), .B2(new_n542), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n425), .A2(new_n435), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n379), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n621), .A2(new_n623), .A3(new_n377), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n598), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n283), .A2(new_n266), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n628), .A2(G472), .B1(new_n285), .B2(new_n283), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n571), .A2(new_n575), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n632), .A2(new_n266), .A3(new_n548), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n583), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n437), .A2(new_n546), .A3(new_n629), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT37), .B(G110), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT94), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(G12));
  AND3_X1   g453(.A1(new_n288), .A2(new_n369), .A3(new_n635), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n618), .A2(new_n620), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n599), .B1(new_n425), .B2(new_n435), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n370), .A2(G900), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(G902), .A3(new_n372), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT95), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT95), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n373), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(KEYINPUT96), .A3(new_n642), .A4(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n642), .A2(new_n618), .A3(new_n620), .A4(new_n647), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n640), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NAND3_X1  g468(.A1(new_n262), .A2(new_n263), .A3(new_n192), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n273), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(KEYINPUT98), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(KEYINPUT98), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G472), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n589), .A2(KEYINPUT32), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n647), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n369), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n622), .B(KEYINPUT38), .Z(new_n669));
  NOR3_X1   g483(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n543), .A2(new_n379), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n494), .B2(new_n499), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n634), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n670), .B(new_n674), .C1(KEYINPUT40), .C2(new_n667), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  AND3_X1   g490(.A1(new_n487), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT88), .B1(new_n487), .B2(KEYINPUT20), .ZN(new_n678));
  INV_X1    g492(.A(new_n493), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n611), .B(new_n647), .C1(new_n680), .C2(new_n619), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n623), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n640), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  OR2_X1    g498(.A1(new_n367), .A2(new_n361), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n367), .A2(new_n361), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n685), .A2(new_n290), .A3(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n612), .A2(new_n288), .A3(new_n586), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n624), .A2(new_n288), .A3(new_n586), .A4(new_n687), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR2_X1   g506(.A1(new_n545), .A2(new_n377), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n685), .A2(new_n290), .A3(new_n686), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n623), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n288), .A3(new_n635), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n581), .A2(new_n582), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n547), .ZN(new_n700));
  INV_X1    g514(.A(new_n585), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n583), .A2(KEYINPUT101), .A3(new_n585), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n264), .A2(new_n257), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n192), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n274), .A2(new_n282), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n285), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT100), .B(G472), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n283), .B2(new_n266), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n704), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n694), .A2(new_n377), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n622), .A3(new_n672), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n628), .A2(new_n710), .B1(new_n285), .B2(new_n707), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n642), .A3(new_n687), .A4(new_n635), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n719), .B2(new_n681), .ZN(new_n720));
  INV_X1    g534(.A(new_n647), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n610), .B(new_n721), .C1(new_n494), .C2(new_n499), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n709), .A2(new_n712), .A3(new_n634), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT102), .A4(new_n695), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NOR2_X1   g540(.A1(new_n344), .A2(new_n355), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n368), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n425), .A2(new_n435), .A3(new_n379), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n729), .A2(new_n291), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n288), .A2(new_n722), .A3(new_n731), .A4(new_n586), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n601), .A2(KEYINPUT42), .A3(new_n611), .A4(new_n647), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n425), .A2(new_n435), .A3(new_n379), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n368), .A2(new_n728), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n290), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n271), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n265), .A2(new_n266), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n255), .B1(new_n279), .B2(new_n250), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n258), .B1(new_n741), .B2(new_n192), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n742), .B2(KEYINPUT29), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n270), .B1(new_n743), .B2(G472), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n704), .B1(new_n745), .B2(new_n663), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n732), .A2(new_n733), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n209), .ZN(G33));
  NOR2_X1   g562(.A1(new_n621), .A2(new_n721), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n288), .A2(new_n749), .A3(new_n731), .A4(new_n586), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  INV_X1    g565(.A(new_n362), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n727), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n356), .B2(new_n359), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n686), .B1(new_n756), .B2(new_n758), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n290), .A4(new_n666), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n680), .A2(new_n619), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n611), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n601), .A2(KEYINPUT43), .A3(new_n610), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n629), .A2(new_n634), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(KEYINPUT44), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n730), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n666), .A2(new_n290), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT105), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n764), .A2(new_n771), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  OR3_X1    g593(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n291), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT47), .B1(new_n775), .B2(new_n291), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n288), .A2(new_n681), .A3(new_n586), .A4(new_n730), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NAND2_X1  g598(.A1(new_n685), .A2(new_n686), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT49), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT49), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n380), .A2(new_n290), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n786), .A2(new_n787), .A3(new_n704), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n766), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n665), .A3(new_n669), .A4(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n640), .B1(new_n652), .B2(new_n682), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n672), .A2(new_n622), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n634), .A2(new_n647), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT108), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n729), .A2(new_n291), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n664), .A2(new_n793), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n725), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n688), .A2(new_n691), .A3(new_n696), .A4(new_n715), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n747), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n494), .A2(new_n499), .A3(new_n543), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n601), .A2(new_n611), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n494), .A2(KEYINPUT106), .A3(new_n499), .A4(new_n543), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n436), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n595), .A2(new_n597), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n587), .A3(new_n636), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n499), .A2(new_n647), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n634), .A2(new_n543), .A3(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n369), .A2(new_n814), .A3(new_n735), .A4(new_n618), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n288), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n722), .A2(new_n723), .A3(new_n731), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n750), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT107), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n802), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n800), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n801), .A2(new_n747), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n587), .A2(new_n636), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n629), .A2(new_n586), .A3(new_n369), .A4(new_n436), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n803), .A2(new_n804), .B1(new_n601), .B2(new_n611), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(new_n807), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n818), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT110), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n812), .A2(new_n837), .A3(new_n818), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n829), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n798), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n792), .A2(new_n725), .A3(new_n799), .A4(new_n797), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n828), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n688), .A2(new_n696), .A3(new_n715), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n732), .A2(new_n733), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n738), .A2(new_n746), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT53), .A4(new_n691), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n437), .A2(new_n546), .ZN(new_n850));
  INV_X1    g664(.A(new_n586), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n745), .B2(new_n663), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n595), .A2(new_n634), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n635), .B(new_n708), .C1(new_n593), .C2(new_n711), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n681), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n856), .A2(new_n731), .B1(new_n815), .B2(new_n288), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n857), .A3(new_n750), .A4(new_n811), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n837), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT110), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n849), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n841), .A2(new_n842), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT111), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n826), .A2(new_n827), .A3(new_n844), .A4(new_n863), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n858), .A2(new_n801), .A3(new_n747), .A4(KEYINPUT107), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n822), .B1(new_n802), .B2(new_n819), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n825), .A3(new_n862), .ZN(new_n868));
  INV_X1    g682(.A(new_n824), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(new_n825), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n864), .B1(new_n870), .B2(new_n827), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n769), .A2(new_n374), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n713), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n669), .A2(new_n599), .A3(new_n687), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT112), .ZN(new_n876));
  OR3_X1    g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n873), .B2(new_n876), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n785), .A2(new_n730), .A3(new_n291), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n665), .A2(new_n586), .A3(new_n374), .A4(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n601), .A3(new_n611), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n872), .A2(new_n880), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n855), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n872), .A2(KEYINPUT113), .A3(new_n723), .A4(new_n880), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n873), .A2(new_n730), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n780), .A2(new_n781), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n785), .A2(new_n290), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n879), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n872), .A2(new_n746), .A3(new_n880), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT48), .Z(new_n896));
  INV_X1    g710(.A(new_n695), .ZN(new_n897));
  OAI221_X1 g711(.A(new_n371), .B1(new_n806), .B2(new_n881), .C1(new_n873), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n892), .B2(new_n893), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n871), .A2(new_n894), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n791), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NAND3_X1  g717(.A1(new_n826), .A2(new_n844), .A3(new_n863), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(G210), .A3(G902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n434), .B(new_n388), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n370), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n863), .A2(new_n844), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT53), .B1(new_n867), .B2(new_n800), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n864), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n362), .B(KEYINPUT57), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n365), .A2(new_n366), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n863), .A2(new_n844), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n266), .B1(new_n921), .B2(new_n826), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n754), .A2(new_n755), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n911), .B1(new_n920), .B2(new_n924), .ZN(G54));
  NAND2_X1  g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT114), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n904), .A2(G902), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n616), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT115), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n911), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n922), .A2(new_n932), .A3(new_n616), .A4(new_n927), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(G60));
  INV_X1    g748(.A(new_n606), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n609), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n871), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n937), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n915), .B2(new_n864), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n911), .A3(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT118), .ZN(new_n943));
  XOR2_X1   g757(.A(KEYINPUT117), .B(KEYINPUT60), .Z(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(new_n944), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n904), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n911), .B1(new_n946), .B2(new_n584), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n632), .B(KEYINPUT119), .Z(new_n948));
  OAI211_X1 g762(.A(new_n945), .B(new_n948), .C1(new_n913), .C2(new_n914), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n911), .ZN(new_n951));
  INV_X1    g765(.A(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n921), .B2(new_n826), .ZN(new_n953));
  INV_X1    g767(.A(new_n584), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n951), .B(new_n949), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n376), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n801), .A2(new_n812), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT120), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n434), .B1(G898), .B2(new_n370), .ZN(new_n965));
  XNOR2_X1  g779(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n964), .B(new_n967), .ZN(G69));
  NAND2_X1  g782(.A1(new_n240), .A2(new_n241), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n469), .A2(new_n470), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n667), .A2(new_n730), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n852), .A2(new_n808), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n778), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n778), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n783), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n792), .A2(KEYINPUT123), .A3(new_n725), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT123), .B1(new_n792), .B2(new_n725), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n675), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(KEYINPUT62), .A3(new_n675), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n977), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n971), .B1(new_n985), .B2(G953), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n848), .A2(new_n750), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n778), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n764), .A2(new_n793), .A3(new_n746), .A4(new_n777), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n988), .A2(new_n783), .A3(new_n980), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n643), .B1(new_n990), .B2(new_n370), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(new_n971), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n643), .B1(new_n339), .B2(G953), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n986), .A2(new_n992), .A3(KEYINPUT125), .A4(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n971), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n983), .A2(new_n984), .ZN(new_n997));
  INV_X1    g811(.A(new_n976), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n778), .A2(new_n972), .A3(new_n974), .ZN(new_n999));
  AOI22_X1  g813(.A1(new_n998), .A2(new_n999), .B1(new_n889), .B2(new_n782), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n996), .B1(new_n1001), .B2(new_n370), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT125), .B1(new_n991), .B2(new_n971), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n993), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n995), .A2(new_n1004), .ZN(G72));
  INV_X1    g819(.A(new_n252), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n741), .A2(new_n192), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n868), .B(new_n1011), .C1(new_n869), .C2(new_n825), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n989), .A2(new_n783), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n963), .A2(new_n980), .A3(new_n988), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(KEYINPUT127), .A3(new_n1009), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1006), .ZN(new_n1016));
  AOI21_X1  g830(.A(KEYINPUT127), .B1(new_n1014), .B2(new_n1009), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n951), .B(new_n1012), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT126), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1010), .B1(new_n985), .B2(new_n963), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1007), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1009), .B1(new_n1001), .B2(new_n962), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1023), .A2(KEYINPUT126), .A3(new_n1007), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1018), .B1(new_n1022), .B2(new_n1024), .ZN(G57));
endmodule


