//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G20), .A3(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n223), .B(new_n227), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n220), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT69), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(G1), .C2(new_n204), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G58), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT70), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT70), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n204), .A2(G33), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR3_X1   g0067(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n265), .A2(new_n267), .B1(new_n268), .B2(new_n204), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n253), .A2(new_n254), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n256), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G222), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G223), .A3(G1698), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n275), .B(new_n276), .C1(new_n210), .C2(new_n273), .ZN(new_n277));
  AND2_X1   g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n254), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n203), .A2(new_n286), .B1(new_n226), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n283), .B1(G226), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n272), .A2(KEYINPUT9), .B1(G200), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n280), .A2(G190), .A3(new_n289), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n291), .B(new_n292), .C1(KEYINPUT9), .C2(new_n272), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n272), .B1(new_n297), .B2(new_n290), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G179), .B2(new_n290), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n249), .A2(KEYINPUT72), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT72), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n302), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n271), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(G68), .C1(G1), .C2(new_n204), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n208), .A2(G20), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n306), .B1(new_n263), .B2(new_n210), .C1(new_n267), .C2(new_n251), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT11), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n307), .A2(new_n308), .A3(new_n271), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n307), .B2(new_n271), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n203), .A2(G13), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n312), .A2(new_n306), .A3(KEYINPUT12), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n301), .A2(new_n303), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n208), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n313), .B1(new_n315), .B2(KEYINPUT12), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n226), .A2(new_n287), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n282), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n321), .A3(new_n282), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(G238), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  OAI211_X1 g0125(.A(G232), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(G226), .B(new_n274), .C1(new_n324), .C2(new_n325), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n279), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n281), .B1(new_n226), .B2(new_n287), .ZN(new_n331));
  INV_X1    g0131(.A(new_n282), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n323), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n209), .B1(new_n288), .B2(new_n321), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n283), .B1(new_n336), .B2(new_n320), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n330), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n317), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G200), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n335), .B2(new_n339), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n317), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  AND4_X1   g0148(.A1(new_n338), .A2(new_n323), .A3(new_n330), .A4(new_n333), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n338), .B1(new_n337), .B2(new_n330), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(G169), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n335), .A2(new_n339), .A3(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n348), .B1(new_n340), .B2(G169), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  OAI211_X1 g0157(.A(G223), .B(new_n274), .C1(new_n324), .C2(new_n325), .ZN(new_n358));
  OAI211_X1 g0158(.A(G226), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G87), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n279), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n288), .A2(G232), .B1(new_n331), .B2(new_n332), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n362), .A2(G190), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n343), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n357), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(G190), .A3(new_n363), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n333), .B1(new_n231), .B2(new_n319), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n279), .B2(new_n361), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(KEYINPUT75), .C1(new_n369), .C2(new_n343), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n259), .A2(G58), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT70), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(new_n376), .A3(new_n255), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n250), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT74), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n249), .B1(new_n261), .B2(new_n262), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(new_n376), .A3(new_n255), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n271), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n324), .A2(new_n325), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n386), .B2(new_n204), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g0188(.A(G33), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT3), .A2(G33), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n257), .A2(new_n208), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n266), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n385), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n384), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n371), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G179), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n362), .A2(new_n409), .A3(new_n363), .ZN(new_n410));
  AOI21_X1  g0210(.A(G169), .B1(new_n362), .B2(new_n363), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT18), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n390), .A2(new_n204), .A3(new_n391), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n208), .B1(new_n416), .B2(new_n392), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n402), .B1(new_n417), .B2(new_n399), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n404), .A3(new_n271), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n380), .A2(new_n382), .A3(new_n381), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n382), .B1(new_n380), .B2(new_n381), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n410), .A2(new_n411), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n405), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n408), .A2(new_n413), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n273), .A2(G232), .A3(new_n274), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n273), .A2(G238), .A3(G1698), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n386), .A2(G107), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n279), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n333), .B1(new_n211), .B2(new_n319), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G200), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n304), .B(G77), .C1(G1), .C2(new_n204), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT8), .B(G58), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n444), .A2(new_n263), .B1(new_n204), .B2(new_n210), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n271), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n314), .A2(new_n210), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n438), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n434), .B1(new_n279), .B2(new_n432), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G190), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n437), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n433), .A2(new_n435), .A3(new_n409), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n448), .C1(G169), .C2(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n300), .A2(new_n356), .A3(new_n428), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n250), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n203), .A2(G33), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n249), .A2(new_n460), .A3(new_n254), .A4(new_n253), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(new_n458), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT76), .ZN(new_n464));
  OAI21_X1  g0264(.A(G107), .B1(new_n387), .B2(new_n393), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n267), .A2(new_n210), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT6), .ZN(new_n467));
  AND2_X1   g0267(.A1(G97), .A2(G107), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G97), .A2(G107), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n466), .B1(new_n473), .B2(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n464), .B1(new_n475), .B2(new_n271), .ZN(new_n476));
  AOI211_X1 g0276(.A(KEYINPUT76), .B(new_n385), .C1(new_n465), .C2(new_n474), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n203), .A2(G45), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(new_n318), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n482), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n331), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G244), .B(new_n274), .C1(new_n324), .C2(new_n325), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n274), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  AOI211_X1 g0294(.A(G190), .B(new_n487), .C1(new_n279), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n279), .ZN(new_n496));
  INV_X1    g0296(.A(new_n487), .ZN(new_n497));
  AOI21_X1  g0297(.A(G200), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n478), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n466), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n471), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  XNOR2_X1  g0302(.A(G97), .B(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n467), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n501), .B1(new_n504), .B2(new_n204), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n471), .B1(new_n416), .B2(new_n392), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n271), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n475), .A2(new_n464), .A3(new_n271), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n462), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n496), .A2(new_n409), .A3(new_n497), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n487), .B1(new_n494), .B2(new_n279), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(G169), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n457), .B1(new_n500), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n509), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n463), .C1(new_n495), .C2(new_n498), .ZN(new_n517));
  AOI211_X1 g0317(.A(G179), .B(new_n487), .C1(new_n279), .C2(new_n494), .ZN(new_n518));
  AOI21_X1  g0318(.A(G169), .B1(new_n496), .B2(new_n497), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n478), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n521), .A3(KEYINPUT77), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n204), .B1(new_n328), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n469), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n204), .B(G68), .C1(new_n324), .C2(new_n325), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n523), .B1(new_n263), .B2(new_n458), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n271), .B1(new_n314), .B2(new_n444), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n249), .A2(new_n460), .ZN(new_n532));
  INV_X1    g0332(.A(new_n444), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT78), .A4(new_n385), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT78), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n461), .B2(new_n444), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT79), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n531), .A2(KEYINPUT79), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G244), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n542));
  OAI211_X1 g0342(.A(G238), .B(new_n274), .C1(new_n324), .C2(new_n325), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n279), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n279), .A2(new_n484), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G250), .B1(new_n331), .B2(new_n484), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(G179), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n297), .B2(new_n549), .ZN(new_n551));
  INV_X1    g0351(.A(new_n549), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G190), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n343), .B1(new_n546), .B2(new_n548), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n530), .A2(new_n271), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n314), .A2(new_n444), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n532), .A2(G87), .A3(new_n385), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n541), .A2(new_n551), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n515), .A2(new_n522), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G270), .B(new_n318), .C1(new_n481), .C2(new_n482), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n562), .A2(new_n486), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n274), .C1(new_n324), .C2(new_n325), .ZN(new_n564));
  OAI211_X1 g0364(.A(G264), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n565));
  INV_X1    g0365(.A(G303), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n273), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n279), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n297), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n492), .B(new_n204), .C1(G33), .C2(new_n458), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT80), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT20), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(G20), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n574), .A3(new_n271), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n571), .B2(new_n572), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n571), .A2(new_n572), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n570), .A2(new_n574), .A3(new_n271), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n203), .B2(G33), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n573), .A2(new_n314), .B1(new_n304), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n579), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n569), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n563), .A2(new_n568), .A3(G179), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n583), .B2(new_n584), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n569), .B(KEYINPUT21), .C1(new_n583), .C2(new_n584), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n204), .B(G87), .C1(new_n324), .C2(new_n325), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g0395(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n596), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n594), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n204), .B2(G107), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n471), .A2(KEYINPUT23), .A3(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G20), .B2(new_n544), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n593), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g0407(.A(KEYINPUT24), .B(new_n605), .C1(new_n597), .C2(new_n599), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n271), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n461), .A2(new_n471), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT25), .B1(new_n250), .B2(new_n471), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT84), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI211_X1 g0413(.A(KEYINPUT84), .B(KEYINPUT25), .C1(new_n250), .C2(new_n471), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n471), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n617), .B(KEYINPUT83), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n610), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(G264), .B(new_n318), .C1(new_n481), .C2(new_n482), .ZN(new_n621));
  NOR2_X1   g0421(.A1(G250), .A2(G1698), .ZN(new_n622));
  INV_X1    g0422(.A(G257), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n623), .B2(G1698), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n273), .B1(G33), .B2(G294), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n486), .B(new_n621), .C1(new_n625), .C2(new_n318), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n343), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G190), .B2(new_n626), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n609), .A2(new_n620), .A3(new_n628), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n615), .A2(new_n618), .B1(new_n471), .B2(new_n461), .ZN(new_n630));
  INV_X1    g0430(.A(new_n599), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n598), .A2(new_n594), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n606), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT24), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n600), .A2(new_n593), .A3(new_n606), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n630), .B1(new_n636), .B2(new_n271), .ZN(new_n637));
  OR3_X1    g0437(.A1(new_n626), .A2(KEYINPUT85), .A3(new_n409), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n626), .A2(G169), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT85), .B1(new_n626), .B2(new_n409), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n629), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n583), .A2(new_n584), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n563), .A2(new_n568), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n645), .B(new_n647), .C1(new_n341), .C2(new_n646), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n592), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n456), .A2(new_n561), .A3(new_n650), .ZN(G372));
  NAND2_X1  g0451(.A1(new_n552), .A2(new_n409), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n549), .A2(new_n297), .ZN(new_n653));
  INV_X1    g0453(.A(new_n540), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n538), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n639), .B(KEYINPUT85), .C1(new_n409), .C2(new_n626), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n385), .B1(new_n634), .B2(new_n635), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n638), .B(new_n656), .C1(new_n657), .C2(new_n630), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(new_n587), .A3(new_n590), .A4(new_n591), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n549), .A2(G200), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n531), .A4(new_n557), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT86), .B1(new_n554), .B2(new_n558), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n553), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n517), .A2(new_n521), .A3(new_n629), .A4(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n655), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n559), .A2(new_n553), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n655), .A2(new_n478), .A3(new_n520), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT87), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n655), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n672), .B2(new_n521), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT87), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n560), .A2(new_n514), .A3(new_n674), .A4(KEYINPUT26), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n456), .B1(new_n667), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n299), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT88), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n413), .A2(KEYINPUT88), .A3(new_n426), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n454), .ZN(new_n685));
  OAI21_X1  g0485(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT14), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n352), .A3(new_n351), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n346), .A2(new_n685), .B1(new_n688), .B2(new_n347), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n405), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT17), .B1(new_n371), .B2(new_n405), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n684), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n694), .A2(new_n695), .B1(new_n295), .B2(new_n294), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n678), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n677), .A2(new_n698), .ZN(G369));
  OR3_X1    g0499(.A1(new_n312), .A2(KEYINPUT27), .A3(G20), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT27), .B1(new_n312), .B2(G20), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(G213), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OR3_X1    g0505(.A1(new_n592), .A2(new_n645), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n592), .A2(new_n648), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n645), .A2(new_n705), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g0509(.A(KEYINPUT90), .B(G330), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n637), .A2(new_n705), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n644), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n715), .A2(new_n716), .B1(new_n658), .B2(new_n705), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n592), .A2(new_n704), .ZN(new_n720));
  INV_X1    g0520(.A(new_n658), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n705), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n221), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G41), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n526), .A2(G116), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G1), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n224), .B2(new_n726), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  INV_X1    g0530(.A(new_n655), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n521), .A2(new_n517), .A3(new_n629), .A4(new_n665), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n659), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n704), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n588), .A2(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n623), .A2(G1698), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G250), .B2(G1698), .ZN(new_n740));
  INV_X1    g0540(.A(G294), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n386), .B1(new_n389), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n279), .ZN(new_n743));
  AND4_X1   g0543(.A1(new_n546), .A2(new_n548), .A3(new_n743), .A4(new_n621), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT92), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n563), .A2(new_n568), .A3(new_n745), .A4(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n738), .A2(new_n512), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n738), .A2(new_n746), .A3(new_n744), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n646), .A2(new_n549), .A3(new_n409), .A4(new_n626), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n512), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n704), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(KEYINPUT31), .B(new_n704), .C1(new_n749), .C2(new_n753), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n515), .A2(new_n522), .A3(new_n560), .A4(new_n705), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n649), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n710), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n672), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(KEYINPUT26), .A3(new_n514), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n669), .A2(KEYINPUT93), .A3(new_n670), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT93), .B1(new_n669), .B2(new_n670), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n733), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n736), .B1(new_n767), .B2(new_n705), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n737), .A2(new_n761), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n730), .B1(new_n769), .B2(G1), .ZN(G364));
  INV_X1    g0570(.A(G13), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n771), .A2(new_n285), .A3(G20), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n773), .A2(G1), .A3(new_n774), .ZN(new_n775));
  OR3_X1    g0575(.A1(new_n725), .A2(new_n775), .A3(KEYINPUT95), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT95), .B1(new_n725), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(G355), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(G355), .A2(new_n780), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n221), .A2(new_n273), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G116), .B2(new_n221), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n247), .A2(G45), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n724), .A2(new_n273), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n285), .B2(new_n225), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n297), .A2(KEYINPUT98), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n204), .B1(KEYINPUT98), .B2(new_n297), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n254), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n779), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G179), .A2(G200), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT100), .ZN(new_n803));
  OAI21_X1  g0603(.A(G20), .B1(new_n803), .B2(new_n341), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT101), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT102), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT102), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G97), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n803), .A2(new_n204), .A3(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n204), .A2(new_n409), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(G190), .A3(G200), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT99), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(KEYINPUT99), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n814), .B1(new_n251), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n815), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n822), .A2(G190), .A3(G200), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n341), .A3(G200), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n273), .B1(new_n824), .B2(new_n210), .C1(new_n257), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n204), .A2(G179), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(G190), .A3(G200), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G87), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n341), .A3(G200), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n822), .A2(G190), .A3(new_n343), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n831), .B1(new_n471), .B2(new_n832), .C1(new_n834), .C2(new_n208), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n812), .A2(KEYINPUT32), .A3(new_n813), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n821), .A2(new_n827), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n810), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT103), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n825), .A2(G322), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n386), .C1(new_n824), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(KEYINPUT33), .A2(G317), .ZN(new_n843));
  AND2_X1   g0643(.A1(KEYINPUT33), .A2(G317), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n833), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G283), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n832), .C1(new_n566), .C2(new_n829), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n842), .B(new_n847), .C1(G329), .C2(new_n811), .ZN(new_n848));
  INV_X1    g0648(.A(new_n805), .ZN(new_n849));
  INV_X1    g0649(.A(G326), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n741), .B2(new_n849), .C1(new_n850), .C2(new_n820), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT104), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n798), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n839), .A2(KEYINPUT104), .A3(new_n851), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n801), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n709), .B2(new_n793), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n711), .A2(new_n779), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n710), .B2(new_n709), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G396));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n791), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n779), .B1(G77), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT105), .Z(new_n864));
  NAND2_X1  g0664(.A1(new_n448), .A2(new_n704), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n452), .A2(new_n454), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT107), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT107), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n685), .A2(new_n704), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n832), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n830), .A2(G107), .B1(new_n873), .B2(G87), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n846), .B2(new_n834), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n273), .B1(new_n823), .B2(G116), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n876), .B1(new_n741), .B2(new_n826), .C1(new_n812), .C2(new_n841), .ZN(new_n877));
  INV_X1    g0677(.A(new_n820), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n875), .B(new_n877), .C1(G303), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n810), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n882));
  AOI22_X1  g0682(.A1(G143), .A2(new_n825), .B1(new_n823), .B2(G159), .ZN(new_n883));
  INV_X1    g0683(.A(G137), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n883), .B1(new_n265), .B2(new_n834), .C1(new_n820), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n886), .A2(KEYINPUT34), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(KEYINPUT34), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n873), .A2(G68), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n273), .C1(new_n251), .C2(new_n829), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G132), .B2(new_n811), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n805), .A2(G58), .ZN(new_n892));
  AND4_X1   g0692(.A1(new_n887), .A2(new_n888), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n881), .A2(new_n882), .A3(new_n893), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n864), .B1(new_n791), .B2(new_n872), .C1(new_n894), .C2(new_n853), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n735), .A2(new_n872), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n868), .A2(new_n869), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n705), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n733), .B2(new_n734), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n760), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n778), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n896), .A2(new_n760), .A3(new_n899), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n895), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT108), .ZN(G384));
  NAND2_X1  g0704(.A1(new_n347), .A2(new_n704), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n346), .A2(new_n355), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n347), .B(new_n704), .C1(new_n688), .C2(new_n345), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n871), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n758), .A2(new_n649), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n756), .A2(new_n757), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT113), .ZN(new_n912));
  INV_X1    g0712(.A(new_n702), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n423), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n428), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n423), .A2(new_n425), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n702), .B(KEYINPUT111), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n423), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n406), .A2(new_n917), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n406), .A2(new_n918), .A3(new_n914), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n917), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n680), .A2(new_n681), .A3(new_n679), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT88), .B1(new_n413), .B2(new_n426), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n692), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n920), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n406), .A2(new_n918), .A3(new_n920), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT37), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n927), .A2(new_n928), .B1(new_n921), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n924), .B1(new_n931), .B2(KEYINPUT38), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT113), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n759), .A2(new_n933), .A3(new_n908), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT114), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n759), .A2(new_n933), .A3(new_n908), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n933), .B1(new_n759), .B2(new_n908), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT38), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n920), .B1(new_n684), .B2(new_n692), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n930), .A2(new_n921), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n945), .B2(new_n924), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(KEYINPUT114), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n916), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT38), .B1(new_n916), .B2(new_n923), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n941), .B1(new_n951), .B2(new_n911), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n456), .A2(new_n759), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n710), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n906), .A2(new_n907), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n898), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n676), .B2(new_n667), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT110), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n454), .A2(new_n704), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT110), .B1(new_n899), .B2(new_n962), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n951), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n684), .A2(new_n919), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n688), .A2(new_n347), .A3(new_n705), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT39), .B1(new_n949), .B2(new_n950), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT39), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n924), .C1(new_n931), .C2(KEYINPUT38), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT112), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(new_n973), .B2(new_n975), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n970), .B1(new_n972), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n456), .B1(new_n737), .B2(new_n768), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n698), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n980), .B(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n956), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n956), .A2(new_n983), .ZN(new_n985));
  OAI21_X1  g0785(.A(G1), .B1(new_n771), .B2(G20), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n473), .A2(KEYINPUT35), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n254), .A2(new_n204), .A3(new_n573), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n473), .B2(KEYINPUT35), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT36), .Z(new_n994));
  NOR3_X1   g0794(.A1(new_n395), .A2(new_n224), .A3(new_n210), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n208), .A2(G50), .ZN(new_n996));
  OAI211_X1 g0796(.A(G1), .B(new_n771), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n987), .A2(new_n994), .A3(new_n997), .ZN(G367));
  NOR2_X1   g0798(.A1(new_n500), .A2(new_n514), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n478), .A2(new_n704), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n514), .A2(new_n704), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n719), .A2(new_n720), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n999), .A2(new_n721), .A3(new_n1000), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n704), .B1(new_n1006), .B2(new_n521), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n1004), .B2(KEYINPUT42), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n558), .A2(new_n704), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n762), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n655), .A2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1005), .A2(new_n1008), .B1(KEYINPUT43), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1013), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1003), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n718), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1017), .B(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n725), .B(KEYINPUT41), .Z(new_n1021));
  NAND3_X1  g0821(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT45), .B1(new_n722), .B2(new_n1003), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n719), .A2(new_n720), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n721), .A2(new_n705), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT44), .B1(new_n1027), .B2(new_n1018), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT44), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n722), .A2(new_n1029), .A3(new_n1003), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1023), .A2(new_n1024), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n718), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n718), .B1(new_n1028), .B2(new_n1030), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1025), .B1(new_n717), .B2(new_n720), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n711), .B(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n769), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1021), .B1(new_n1037), .B2(new_n769), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1020), .B1(new_n1038), .B2(new_n775), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n799), .B1(new_n221), .B2(new_n444), .C1(new_n237), .C2(new_n787), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(new_n779), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n809), .A2(G68), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n273), .B1(new_n824), .B2(new_n251), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G150), .B2(new_n825), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n878), .A2(G143), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n833), .A2(G159), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n873), .A2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n811), .A2(G137), .B1(G58), .B2(new_n830), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1048), .B1(KEYINPUT116), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1042), .B(new_n1050), .C1(KEYINPUT116), .C2(new_n1049), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT46), .B1(new_n830), .B2(G116), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G283), .A2(new_n823), .B1(new_n825), .B2(G303), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n830), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n741), .C2(new_n834), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1052), .B(new_n1055), .C1(G311), .C2(new_n878), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n832), .A2(new_n458), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n273), .B(new_n1057), .C1(new_n811), .C2(G317), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT115), .Z(new_n1059));
  OAI211_X1 g0859(.A(new_n1056), .B(new_n1059), .C1(new_n471), .C2(new_n849), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT47), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n1041), .B1(new_n793), .B2(new_n1012), .C1(new_n1062), .C2(new_n853), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1039), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT117), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1039), .A2(new_n1067), .A3(new_n1063), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1066), .A2(new_n1069), .ZN(G387));
  INV_X1    g0870(.A(new_n727), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n221), .A3(new_n273), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(G107), .B2(new_n221), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT118), .Z(new_n1074));
  OR2_X1    g0874(.A1(new_n234), .A2(new_n285), .ZN(new_n1075));
  AOI211_X1 g0875(.A(G45), .B(new_n1071), .C1(G68), .C2(G77), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n439), .A2(G50), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n787), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1074), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n779), .B1(new_n1080), .B2(new_n800), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n809), .A2(new_n533), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n878), .A2(G159), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n273), .B1(new_n824), .B2(new_n208), .C1(new_n251), .C2(new_n826), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1057), .B(new_n1084), .C1(G77), .C2(new_n830), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT119), .B(G150), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n261), .A2(new_n262), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n811), .A2(new_n1086), .B1(new_n1087), .B2(new_n833), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G303), .A2(new_n823), .B1(new_n825), .B2(G317), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n841), .B2(new_n834), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G322), .B2(new_n878), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT48), .Z(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n846), .B2(new_n849), .C1(new_n741), .C2(new_n829), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT49), .Z(new_n1095));
  OAI221_X1 g0895(.A(new_n386), .B1(new_n832), .B2(new_n573), .C1(new_n812), .C2(new_n850), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1081), .B1(new_n1097), .B2(new_n798), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n717), .A2(new_n793), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1098), .A2(new_n1099), .B1(new_n775), .B2(new_n1036), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1036), .A2(new_n769), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n725), .B(KEYINPUT120), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(KEYINPUT121), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n769), .B2(new_n1036), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT121), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(G393));
  NAND2_X1  g0906(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1018), .A2(new_n794), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n799), .B1(new_n458), .B2(new_n221), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n242), .B2(new_n786), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n808), .A2(new_n210), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n273), .B1(new_n824), .B2(new_n439), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n834), .A2(new_n251), .B1(new_n208), .B2(new_n829), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(G87), .C2(new_n873), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n820), .A2(new_n265), .B1(new_n813), .B2(new_n826), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT51), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n811), .A2(G143), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n834), .A2(new_n566), .B1(new_n846), .B2(new_n829), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n386), .B1(new_n471), .B2(new_n832), .C1(new_n824), .C2(new_n741), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G322), .C2(new_n811), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n573), .B2(new_n849), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n878), .A2(G317), .B1(G311), .B2(new_n825), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT52), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1112), .A2(new_n1121), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n778), .B(new_n1111), .C1(new_n1128), .C2(new_n798), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1108), .A2(new_n775), .B1(new_n1109), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1107), .A2(new_n1101), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n1037), .A3(new_n1102), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(G390));
  AOI21_X1  g0933(.A(new_n962), .B1(new_n767), .B2(new_n959), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n958), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n932), .A2(new_n971), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n761), .A2(new_n872), .A3(new_n957), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n966), .A2(new_n972), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(new_n1139), .C1(new_n979), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n973), .A2(new_n975), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT112), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n964), .A2(new_n965), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n957), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n971), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1137), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n759), .A2(G330), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(new_n908), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1141), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n456), .A2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n981), .A2(new_n698), .A3(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1150), .A2(new_n872), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1134), .B(new_n1139), .C1(new_n1156), .C2(new_n957), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n957), .B1(new_n761), .B2(new_n872), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1146), .B1(new_n1158), .B2(new_n1151), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1155), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1153), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1141), .B(new_n1160), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1102), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1141), .B(new_n775), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n273), .B1(new_n825), .B2(G116), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n831), .A3(new_n889), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n834), .A2(new_n471), .B1(new_n824), .B2(new_n458), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n878), .B2(G283), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT122), .Z(new_n1170));
  AOI211_X1 g0970(.A(new_n1167), .B(new_n1170), .C1(G294), .C2(new_n811), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1112), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n809), .A2(G159), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n830), .A2(new_n1086), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT53), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n824), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n811), .A2(G125), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n386), .B1(new_n825), .B2(G132), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n833), .A2(G137), .B1(G50), .B2(new_n873), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1175), .B(new_n1181), .C1(G128), .C2(new_n878), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1171), .A2(new_n1172), .B1(new_n1173), .B2(new_n1182), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n779), .B1(new_n1087), .B2(new_n862), .C1(new_n1183), .C2(new_n853), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT123), .Z(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n791), .B2(new_n979), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1165), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1164), .A2(new_n1187), .ZN(G378));
  OAI211_X1 g0988(.A(new_n968), .B(new_n969), .C1(new_n1145), .C2(new_n971), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n272), .A2(new_n702), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n296), .A2(new_n299), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n296), .B2(new_n299), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1191), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1196), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n1194), .A3(new_n1190), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n952), .A2(G330), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n937), .C2(new_n947), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1200), .B1(new_n948), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1189), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT114), .B1(new_n940), .B2(new_n946), .ZN(new_n1207));
  AND4_X1   g1007(.A1(KEYINPUT114), .A2(new_n946), .A3(new_n912), .A4(new_n934), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1204), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1201), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n948), .A2(new_n1204), .A3(new_n1200), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n980), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1201), .A2(new_n790), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n779), .B1(G50), .B2(new_n862), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n830), .A2(G77), .B1(new_n873), .B2(G58), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n458), .B2(new_n834), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n386), .A2(new_n284), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n825), .B2(G107), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n444), .B2(new_n824), .C1(new_n812), .C2(new_n846), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1217), .B(new_n1220), .C1(G116), .C2(new_n878), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1042), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G50), .B1(new_n389), .B2(new_n284), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1222), .A2(new_n1223), .B1(new_n1218), .B2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT124), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n829), .A2(new_n1176), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G128), .A2(new_n825), .B1(new_n823), .B2(G137), .ZN(new_n1228));
  INV_X1    g1028(.A(G132), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n834), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1227), .B(new_n1230), .C1(G125), .C2(new_n878), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n808), .B2(new_n265), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n389), .B(new_n284), .C1(new_n832), .C2(new_n813), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n811), .B2(G124), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1226), .B1(new_n1223), .B2(new_n1222), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1215), .B1(new_n1238), .B2(new_n798), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1213), .A2(new_n775), .B1(new_n1214), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1155), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1163), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1102), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1242), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1240), .B1(new_n1244), .B2(new_n1245), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n958), .A2(new_n790), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n779), .B1(G68), .B2(new_n862), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n386), .B1(new_n823), .B2(G150), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n257), .B2(new_n832), .C1(new_n813), .C2(new_n829), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G128), .B2(new_n811), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n808), .B2(new_n251), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT126), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n884), .A2(new_n826), .B1(new_n834), .B2(new_n1176), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G132), .B2(new_n878), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1047), .B1(new_n458), .B2(new_n829), .C1(new_n834), .C2(new_n573), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n273), .B1(new_n823), .B2(G107), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n846), .B2(new_n826), .C1(new_n812), .C2(new_n566), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G294), .C2(new_n878), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1082), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1249), .B1(new_n1263), .B2(new_n798), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1247), .A2(new_n775), .B1(new_n1248), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1247), .B2(new_n1241), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1157), .A2(new_n1159), .A3(KEYINPUT125), .A4(new_n1155), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1021), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1161), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1265), .B1(new_n1269), .B2(new_n1271), .ZN(G381));
  INV_X1    g1072(.A(G390), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G396), .A2(new_n1275), .A3(G393), .A4(G381), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G387), .A2(new_n1276), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n703), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  OAI211_X1 g1082(.A(G378), .B(new_n1240), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1213), .A2(new_n1270), .A3(new_n1242), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1240), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1278), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1279), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1267), .B(new_n1268), .C1(new_n1289), .C2(new_n1160), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1102), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1247), .A2(new_n1241), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1274), .B1(new_n1294), .B2(new_n1265), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1274), .A3(new_n1265), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(G2897), .A3(new_n1280), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1280), .A2(G2897), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1297), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1295), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1065), .A2(new_n1068), .A3(new_n1273), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1065), .A2(KEYINPUT127), .A3(new_n1068), .A4(new_n1273), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(G393), .B(G396), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1039), .A2(G390), .A3(new_n1063), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1064), .B(G390), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1315), .A2(new_n1310), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1300), .A2(new_n1295), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1319), .B1(new_n1288), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1280), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1320), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(KEYINPUT63), .A3(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1304), .A2(new_n1318), .A3(new_n1321), .A4(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1322), .A2(new_n1326), .A3(new_n1323), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1322), .B2(new_n1302), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1327), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1325), .B1(new_n1331), .B2(new_n1318), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1278), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1283), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1323), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1312), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1336), .A2(new_n1320), .A3(new_n1316), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1334), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1314), .A2(new_n1323), .A3(new_n1317), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1320), .B1(new_n1336), .B2(new_n1316), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1283), .A4(new_n1333), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(G402));
endmodule


