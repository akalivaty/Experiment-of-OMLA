

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U552 ( .A(n881), .Z(n519) );
  XNOR2_X1 U553 ( .A(n521), .B(n520), .ZN(n881) );
  NAND2_X1 U554 ( .A1(G8), .A2(n735), .ZN(n810) );
  BUF_X1 U555 ( .A(n545), .Z(n536) );
  XOR2_X1 U556 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  XNOR2_X2 U557 ( .A(n569), .B(KEYINPUT76), .ZN(n974) );
  AND2_X1 U558 ( .A1(n767), .A2(n683), .ZN(n705) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X2 U560 ( .A(KEYINPUT1), .B(n563), .ZN(n573) );
  NOR2_X2 U561 ( .A1(G2104), .A2(n524), .ZN(n532) );
  XNOR2_X1 U562 ( .A(n704), .B(KEYINPUT97), .ZN(n709) );
  NOR2_X1 U563 ( .A1(n974), .A2(n710), .ZN(n717) );
  NOR2_X1 U564 ( .A1(n701), .A2(n700), .ZN(n721) );
  INV_X1 U565 ( .A(KEYINPUT103), .ZN(n733) );
  NOR2_X1 U566 ( .A1(G1966), .A2(n810), .ZN(n744) );
  INV_X1 U567 ( .A(n766), .ZN(n683) );
  OR2_X1 U568 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U569 ( .A1(n881), .A2(G138), .ZN(n523) );
  INV_X1 U570 ( .A(KEYINPUT17), .ZN(n520) );
  XNOR2_X1 U571 ( .A(KEYINPUT66), .B(n559), .ZN(n647) );
  INV_X1 U572 ( .A(KEYINPUT87), .ZN(n531) );
  INV_X1 U573 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G126), .A2(n532), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n529) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U577 ( .A1(G114), .A2(n887), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n524), .A2(G2104), .ZN(n525) );
  XNOR2_X1 U579 ( .A(n525), .B(KEYINPUT67), .ZN(n545) );
  NAND2_X1 U580 ( .A1(G102), .A2(n545), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U583 ( .A(n531), .B(n530), .ZN(n681) );
  BUF_X1 U584 ( .A(n681), .Z(G164) );
  AND2_X1 U585 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U586 ( .A1(n532), .A2(G123), .ZN(n533) );
  XNOR2_X1 U587 ( .A(n533), .B(KEYINPUT18), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G111), .A2(n887), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G135), .A2(n519), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G99), .A2(n536), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n929) );
  XNOR2_X1 U594 ( .A(n929), .B(G2096), .ZN(n541) );
  XNOR2_X1 U595 ( .A(n541), .B(KEYINPUT79), .ZN(n542) );
  OR2_X1 U596 ( .A1(G2100), .A2(n542), .ZN(G156) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  INV_X1 U598 ( .A(G120), .ZN(G236) );
  INV_X1 U599 ( .A(G69), .ZN(G235) );
  INV_X1 U600 ( .A(G108), .ZN(G238) );
  NAND2_X1 U601 ( .A1(G125), .A2(n532), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G113), .A2(n887), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n551) );
  XOR2_X1 U604 ( .A(KEYINPUT68), .B(KEYINPUT23), .Z(n547) );
  NAND2_X1 U605 ( .A1(G101), .A2(n545), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n519), .A2(G137), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n551), .A2(n550), .ZN(G160) );
  NAND2_X1 U610 ( .A1(G7), .A2(G661), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n552), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U612 ( .A(G223), .B(KEYINPUT74), .Z(n833) );
  NAND2_X1 U613 ( .A1(n833), .A2(G567), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n553), .Z(G234) );
  INV_X1 U615 ( .A(G860), .ZN(n606) );
  NOR2_X1 U616 ( .A1(G543), .A2(G651), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT65), .B(n554), .Z(n637) );
  NAND2_X1 U618 ( .A1(n637), .A2(G81), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT12), .ZN(n557) );
  XNOR2_X1 U620 ( .A(KEYINPUT69), .B(G651), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n646), .A2(n561), .ZN(n640) );
  NAND2_X1 U622 ( .A1(G68), .A2(n640), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT13), .ZN(n568) );
  NOR2_X1 U625 ( .A1(G651), .A2(n646), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n647), .A2(G43), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT75), .ZN(n566) );
  NOR2_X1 U628 ( .A1(G543), .A2(n561), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT70), .B(n562), .Z(n563) );
  NAND2_X1 U630 ( .A1(G56), .A2(n573), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U634 ( .A1(n606), .A2(n974), .ZN(G153) );
  NAND2_X1 U635 ( .A1(G90), .A2(n637), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G77), .A2(n640), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT9), .B(n572), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n647), .A2(G52), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(G64), .ZN(n574) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G92), .A2(n637), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G79), .A2(n640), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G54), .A2(n647), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G66), .A2(n573), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n584), .Z(n976) );
  OR2_X1 U652 ( .A1(n976), .A2(G868), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U654 ( .A1(n637), .A2(G89), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT4), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G76), .A2(n640), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT5), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G51), .A2(n647), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G63), .A2(n573), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT6), .B(n593), .Z(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n596), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U665 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U666 ( .A1(n640), .A2(G78), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G53), .A2(n647), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n637), .A2(G91), .ZN(n599) );
  XOR2_X1 U670 ( .A(KEYINPUT72), .B(n599), .Z(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U672 ( .A1(G65), .A2(n573), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(G299) );
  INV_X1 U674 ( .A(G868), .ZN(n662) );
  NOR2_X1 U675 ( .A1(G286), .A2(n662), .ZN(n605) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n607), .A2(n976), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT16), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT77), .B(n609), .Z(G148) );
  NOR2_X1 U682 ( .A1(n974), .A2(G868), .ZN(n610) );
  XNOR2_X1 U683 ( .A(KEYINPUT78), .B(n610), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G868), .A2(n976), .ZN(n611) );
  NOR2_X1 U685 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G559), .A2(n976), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(n974), .ZN(n660) );
  NOR2_X1 U689 ( .A1(G860), .A2(n660), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G80), .A2(n640), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT80), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G55), .A2(n647), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G93), .A2(n637), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G67), .A2(n573), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n663) );
  XOR2_X1 U698 ( .A(n622), .B(n663), .Z(G145) );
  NAND2_X1 U699 ( .A1(G88), .A2(n637), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G75), .A2(n640), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G50), .A2(n647), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G62), .A2(n573), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G166) );
  NAND2_X1 U706 ( .A1(G85), .A2(n637), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G60), .A2(n573), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G47), .A2(n647), .ZN(n631) );
  XNOR2_X1 U710 ( .A(KEYINPUT71), .B(n631), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n640), .A2(G72), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U714 ( .A1(n573), .A2(G61), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT82), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n637), .A2(G86), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G48), .A2(n647), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n640), .A2(G73), .ZN(n641) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U723 ( .A1(n646), .A2(G87), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G49), .A2(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U726 ( .A1(n573), .A2(n650), .ZN(n653) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n651) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(n651), .Z(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(G288) );
  INV_X1 U730 ( .A(G299), .ZN(n720) );
  XNOR2_X1 U731 ( .A(n720), .B(G166), .ZN(n659) );
  XOR2_X1 U732 ( .A(n663), .B(G290), .Z(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(G305), .ZN(n655) );
  XNOR2_X1 U734 ( .A(KEYINPUT83), .B(n655), .ZN(n657) );
  XNOR2_X1 U735 ( .A(G288), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(n899) );
  XOR2_X1 U738 ( .A(n899), .B(n660), .Z(n661) );
  NOR2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n665) );
  NOR2_X1 U740 ( .A1(G868), .A2(n663), .ZN(n664) );
  NOR2_X1 U741 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n667), .ZN(n669) );
  XNOR2_X1 U745 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U747 ( .A1(G2072), .A2(n670), .ZN(G158) );
  XNOR2_X1 U748 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G235), .A2(G236), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT86), .B(n671), .Z(n672) );
  NOR2_X1 U752 ( .A1(G238), .A2(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G57), .A2(n673), .ZN(n837) );
  NAND2_X1 U754 ( .A1(n837), .A2(G567), .ZN(n679) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n675) );
  XNOR2_X1 U756 ( .A(KEYINPUT85), .B(KEYINPUT22), .ZN(n674) );
  XNOR2_X1 U757 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U758 ( .A1(n676), .A2(G218), .ZN(n677) );
  NAND2_X1 U759 ( .A1(G96), .A2(n677), .ZN(n838) );
  NAND2_X1 U760 ( .A1(n838), .A2(G2106), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n839) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U763 ( .A1(n839), .A2(n680), .ZN(n836) );
  NAND2_X1 U764 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G301), .ZN(G171) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  NOR2_X1 U767 ( .A1(n681), .A2(G1384), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n682), .B(KEYINPUT64), .ZN(n767) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n766) );
  INV_X1 U770 ( .A(KEYINPUT93), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n705), .B(n684), .ZN(n712) );
  XNOR2_X1 U772 ( .A(G2078), .B(KEYINPUT25), .ZN(n952) );
  NAND2_X1 U773 ( .A1(n712), .A2(n952), .ZN(n686) );
  INV_X1 U774 ( .A(n705), .ZN(n735) );
  INV_X1 U775 ( .A(G1961), .ZN(n998) );
  NAND2_X1 U776 ( .A1(n735), .A2(n998), .ZN(n685) );
  NAND2_X1 U777 ( .A1(n686), .A2(n685), .ZN(n728) );
  OR2_X1 U778 ( .A1(n728), .A2(G171), .ZN(n687) );
  XNOR2_X1 U779 ( .A(n687), .B(KEYINPUT101), .ZN(n695) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n735), .ZN(n743) );
  NOR2_X1 U781 ( .A1(n744), .A2(n743), .ZN(n689) );
  INV_X1 U782 ( .A(KEYINPUT99), .ZN(n688) );
  XNOR2_X1 U783 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n690), .A2(G8), .ZN(n692) );
  XNOR2_X1 U785 ( .A(KEYINPUT30), .B(KEYINPUT100), .ZN(n691) );
  XNOR2_X1 U786 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n693), .A2(G168), .ZN(n694) );
  NOR2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n697) );
  XOR2_X1 U789 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n696) );
  XNOR2_X1 U790 ( .A(n697), .B(n696), .ZN(n732) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n712), .ZN(n699) );
  XOR2_X1 U792 ( .A(KEYINPUT94), .B(KEYINPUT27), .Z(n698) );
  XOR2_X1 U793 ( .A(n699), .B(n698), .Z(n701) );
  INV_X1 U794 ( .A(G1956), .ZN(n1004) );
  NOR2_X1 U795 ( .A1(n712), .A2(n1004), .ZN(n700) );
  NOR2_X1 U796 ( .A1(n721), .A2(n720), .ZN(n703) );
  XNOR2_X1 U797 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n703), .B(n702), .ZN(n725) );
  AND2_X1 U799 ( .A1(G1341), .A2(n735), .ZN(n704) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n705), .ZN(n707) );
  XNOR2_X1 U801 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n706) );
  XNOR2_X1 U802 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n976), .A2(n717), .ZN(n716) );
  NAND2_X1 U805 ( .A1(G1348), .A2(n735), .ZN(n711) );
  XNOR2_X1 U806 ( .A(n711), .B(KEYINPUT98), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n712), .A2(G2067), .ZN(n713) );
  NAND2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n719) );
  OR2_X1 U810 ( .A1(n976), .A2(n717), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n727) );
  INV_X1 U815 ( .A(KEYINPUT29), .ZN(n726) );
  XNOR2_X1 U816 ( .A(n727), .B(n726), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n728), .A2(G171), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n745) );
  NAND2_X1 U820 ( .A1(G286), .A2(n745), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(n733), .ZN(n740) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n810), .ZN(n737) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U825 ( .A1(G303), .A2(n738), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n741), .A2(G8), .ZN(n742) );
  XNOR2_X1 U828 ( .A(n742), .B(KEYINPUT32), .ZN(n805) );
  NAND2_X1 U829 ( .A1(G8), .A2(n743), .ZN(n748) );
  INV_X1 U830 ( .A(n745), .ZN(n746) );
  NOR2_X1 U831 ( .A1(n744), .A2(n746), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n748), .A2(n747), .ZN(n806) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n979) );
  AND2_X1 U834 ( .A1(n806), .A2(n979), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n805), .A2(n749), .ZN(n753) );
  INV_X1 U836 ( .A(n979), .ZN(n751) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n755), .A2(n750), .ZN(n983) );
  OR2_X1 U840 ( .A1(n751), .A2(n983), .ZN(n752) );
  AND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U842 ( .A(n754), .B(KEYINPUT104), .ZN(n759) );
  NAND2_X1 U843 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  XOR2_X1 U844 ( .A(KEYINPUT105), .B(n756), .Z(n757) );
  NOR2_X1 U845 ( .A1(n810), .A2(n757), .ZN(n760) );
  OR2_X1 U846 ( .A1(n810), .A2(n760), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n763) );
  INV_X1 U848 ( .A(n760), .ZN(n761) );
  AND2_X1 U849 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  XNOR2_X1 U850 ( .A(n764), .B(KEYINPUT106), .ZN(n801) );
  XOR2_X1 U851 ( .A(G1981), .B(KEYINPUT107), .Z(n765) );
  XNOR2_X1 U852 ( .A(G305), .B(n765), .ZN(n972) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U854 ( .A(n768), .B(KEYINPUT88), .ZN(n826) );
  INV_X1 U855 ( .A(n826), .ZN(n795) );
  NAND2_X1 U856 ( .A1(G119), .A2(n532), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G131), .A2(n519), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G107), .A2(n887), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G95), .A2(n536), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n867) );
  NAND2_X1 U863 ( .A1(G1991), .A2(n867), .ZN(n775) );
  XNOR2_X1 U864 ( .A(n775), .B(KEYINPUT91), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G129), .A2(n532), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G117), .A2(n887), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n536), .A2(G105), .ZN(n778) );
  XOR2_X1 U869 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n519), .A2(G141), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n893) );
  AND2_X1 U873 ( .A1(G1996), .A2(n893), .ZN(n783) );
  NOR2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n931) );
  NOR2_X1 U875 ( .A1(n795), .A2(n931), .ZN(n818) );
  INV_X1 U876 ( .A(n818), .ZN(n797) );
  NAND2_X1 U877 ( .A1(n532), .A2(G128), .ZN(n785) );
  XOR2_X1 U878 ( .A(KEYINPUT89), .B(n785), .Z(n787) );
  NAND2_X1 U879 ( .A1(n887), .A2(G116), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U881 ( .A(n788), .B(KEYINPUT35), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G140), .A2(n519), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G104), .A2(n536), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT34), .B(n791), .Z(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n794), .B(KEYINPUT36), .ZN(n896) );
  XOR2_X1 U888 ( .A(G2067), .B(KEYINPUT37), .Z(n823) );
  NAND2_X1 U889 ( .A1(n896), .A2(n823), .ZN(n936) );
  NOR2_X1 U890 ( .A1(n795), .A2(n936), .ZN(n796) );
  XOR2_X1 U891 ( .A(KEYINPUT90), .B(n796), .Z(n821) );
  NAND2_X1 U892 ( .A1(n797), .A2(n821), .ZN(n799) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n985) );
  AND2_X1 U894 ( .A1(n985), .A2(n826), .ZN(n798) );
  OR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n815) );
  NOR2_X1 U896 ( .A1(n972), .A2(n815), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n831) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XOR2_X1 U899 ( .A(n802), .B(KEYINPUT92), .Z(n803) );
  XNOR2_X1 U900 ( .A(KEYINPUT24), .B(n803), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n804), .A2(n810), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U903 ( .A1(G2090), .A2(G303), .ZN(n807) );
  NAND2_X1 U904 ( .A1(G8), .A2(n807), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n811) );
  AND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n829) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n893), .ZN(n925) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n867), .ZN(n933) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U912 ( .A1(n933), .A2(n816), .ZN(n817) );
  NOR2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n925), .A2(n819), .ZN(n820) );
  XNOR2_X1 U915 ( .A(KEYINPUT39), .B(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n825) );
  NOR2_X1 U917 ( .A1(n896), .A2(n823), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT108), .B(n824), .Z(n937) );
  NAND2_X1 U919 ( .A1(n825), .A2(n937), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  AND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U923 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U926 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n839), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n843) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U940 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2078), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1976), .B(G1986), .Z(n849) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n859) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G2474), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1981), .B(KEYINPUT110), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U949 ( .A(G1971), .B(G1956), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U953 ( .A(KEYINPUT112), .B(KEYINPUT111), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U956 ( .A1(n532), .A2(G124), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G112), .A2(n887), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U960 ( .A1(G136), .A2(n519), .ZN(n864) );
  NAND2_X1 U961 ( .A1(G100), .A2(n536), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U963 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n869) );
  XNOR2_X1 U965 ( .A(n867), .B(n929), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n878) );
  NAND2_X1 U967 ( .A1(n536), .A2(G103), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n870), .B(KEYINPUT114), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G139), .A2(n519), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G127), .A2(n532), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G115), .A2(n887), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n920) );
  XOR2_X1 U976 ( .A(n878), .B(n920), .Z(n880) );
  XNOR2_X1 U977 ( .A(G164), .B(G162), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n892) );
  NAND2_X1 U979 ( .A1(G142), .A2(n519), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G106), .A2(n536), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(KEYINPUT45), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G130), .A2(n532), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n890) );
  NAND2_X1 U985 ( .A1(G118), .A2(n887), .ZN(n888) );
  XNOR2_X1 U986 ( .A(KEYINPUT113), .B(n888), .ZN(n889) );
  NOR2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(n892), .B(n891), .Z(n895) );
  XOR2_X1 U989 ( .A(G160), .B(n893), .Z(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U993 ( .A(n899), .B(G286), .Z(n901) );
  XNOR2_X1 U994 ( .A(G171), .B(n976), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n974), .B(n902), .Z(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U998 ( .A(KEYINPUT109), .B(G2446), .Z(n905) );
  XNOR2_X1 U999 ( .A(G2435), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2430), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G2454), .B(G2427), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n908), .B(G2443), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G57), .ZN(G237) );
  INV_X1 U1017 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G2072), .B(n920), .Z(n922) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1021 ( .A(KEYINPUT50), .B(n923), .Z(n942) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n926), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(KEYINPUT115), .ZN(n935) );
  XOR2_X1 U1026 ( .A(G2084), .B(G160), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1033 ( .A(KEYINPUT116), .B(n940), .Z(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n943), .ZN(n944) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n967), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n945), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(G34), .Z(n947) );
  XNOR2_X1 U1040 ( .A(G2084), .B(KEYINPUT54), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(n947), .B(n946), .ZN(n965) );
  XNOR2_X1 U1042 ( .A(G2090), .B(G35), .ZN(n963) );
  XNOR2_X1 U1043 ( .A(G32), .B(G1996), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(n948), .B(KEYINPUT119), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(G28), .A2(n951), .ZN(n955) );
  XOR2_X1 U1049 ( .A(G27), .B(n952), .Z(n953) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(n953), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G25), .B(G1991), .Z(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT117), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n961), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1060 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n970), .ZN(n1027) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XOR2_X1 U1064 ( .A(G1966), .B(G168), .Z(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT57), .B(n973), .Z(n995) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n974), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT123), .ZN(n990) );
  XNOR2_X1 U1069 ( .A(n976), .B(G1348), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n977), .B(KEYINPUT121), .ZN(n988) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G299), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT122), .B(n986), .Z(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G301), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n993), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n1025) );
  XNOR2_X1 U1085 ( .A(G5), .B(n998), .ZN(n1012) );
  XNOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n999), .B(G4), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G6), .B(G1981), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(KEYINPUT126), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1093 ( .A(G20), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G21), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G1986), .B(KEYINPUT127), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(G24), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT61), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G16), .B(KEYINPUT125), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

