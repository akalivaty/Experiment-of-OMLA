//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT16), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n197), .A3(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT78), .A4(G146), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n206), .B(KEYINPUT74), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT24), .B(G110), .Z(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n203), .A2(new_n204), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT75), .B1(new_n205), .B2(G119), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n217), .C1(new_n218), .C2(new_n216), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(KEYINPUT76), .A3(new_n216), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n221), .A3(G110), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(new_n225), .A3(KEYINPUT79), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n215), .B1(new_n208), .B2(G128), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n206), .B1(new_n228), .B2(KEYINPUT23), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n229), .A2(new_n217), .B1(new_n220), .B2(new_n210), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(new_n224), .A3(G110), .A4(new_n222), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n223), .A2(KEYINPUT77), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n203), .A2(new_n204), .A3(new_n212), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n227), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n226), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n193), .A2(new_n195), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n199), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n240));
  INV_X1    g054(.A(G110), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT80), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(KEYINPUT80), .A3(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n211), .B1(new_n207), .B2(new_n210), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n202), .B(new_n239), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n236), .A2(new_n237), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n237), .B1(new_n236), .B2(new_n248), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n191), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G902), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n236), .A2(new_n248), .A3(new_n190), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n252), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT73), .B(G217), .Z(new_n259));
  INV_X1    g073(.A(G234), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G902), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n251), .A2(new_n253), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n262), .A2(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT9), .B(G234), .Z(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n252), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G221), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT82), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G469), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n275));
  INV_X1    g089(.A(G107), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(G104), .ZN(new_n277));
  INV_X1    g091(.A(G104), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(G107), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n279));
  OAI22_X1  g093(.A1(new_n278), .A2(G107), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G101), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n282), .A2(KEYINPUT4), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n284));
  XNOR2_X1  g098(.A(G143), .B(G146), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n199), .A2(G143), .ZN(new_n289));
  INV_X1    g103(.A(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G146), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OR2_X1    g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n292), .A2(new_n284), .A3(new_n286), .A4(new_n293), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G101), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n277), .A2(new_n279), .A3(new_n280), .A4(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(KEYINPUT84), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n282), .A2(KEYINPUT4), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n283), .B(new_n297), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n278), .A2(G107), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n276), .A2(G104), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n285), .A2(new_n307), .A3(G128), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n290), .A2(KEYINPUT1), .A3(G146), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n308), .B(new_n309), .C1(G128), .C2(new_n285), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT84), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n299), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n299), .A2(new_n311), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n306), .B(new_n310), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G128), .B1(new_n289), .B2(new_n291), .ZN(new_n317));
  INV_X1    g131(.A(new_n309), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT67), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n309), .B(new_n320), .C1(new_n285), .C2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n322), .B2(new_n308), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n277), .A2(new_n280), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(KEYINPUT84), .A3(new_n298), .A4(new_n279), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n299), .A2(new_n311), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n305), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT11), .ZN(new_n329));
  INV_X1    g143(.A(G134), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(G137), .ZN(new_n331));
  INV_X1    g145(.A(G137), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT11), .A3(G134), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(G137), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G131), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n331), .A2(new_n333), .A3(new_n338), .A4(new_n334), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(KEYINPUT65), .A3(G131), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n302), .A2(new_n316), .A3(new_n328), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT85), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n315), .A2(new_n314), .B1(new_n323), .B2(new_n327), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n343), .A4(new_n302), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n188), .A2(G227), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n350), .B(new_n351), .Z(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n302), .A2(new_n316), .A3(new_n328), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n354), .A2(new_n355), .A3(new_n342), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n354), .B2(new_n342), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n322), .A2(new_n308), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n314), .B1(new_n327), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n342), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT12), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(KEYINPUT12), .A3(new_n342), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n345), .A2(new_n348), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n353), .A2(new_n358), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT87), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n349), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n352), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n354), .A2(new_n342), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT86), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n354), .A2(new_n355), .A3(new_n342), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n349), .A3(new_n352), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n273), .B1(new_n367), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n352), .B1(new_n375), .B2(new_n349), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n349), .A2(new_n352), .A3(new_n368), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n273), .B(new_n252), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n273), .A2(new_n252), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n272), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n267), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G237), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n188), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n290), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT92), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT18), .A2(G131), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n238), .B(G146), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n392), .B(new_n338), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n203), .A2(new_n204), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(KEYINPUT17), .A3(G131), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(G113), .B(G122), .Z(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT94), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT93), .B(G104), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n398), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n238), .B(KEYINPUT19), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n202), .B1(new_n412), .B2(G146), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n399), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n408), .B1(new_n414), .B2(new_n397), .ZN(new_n415));
  AOI21_X1  g229(.A(G475), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n252), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT20), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n419), .A3(new_n252), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n410), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n409), .B1(new_n398), .B2(new_n404), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n252), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT95), .B(G475), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G116), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT96), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(KEYINPUT68), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G122), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n276), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(G107), .A3(new_n436), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(KEYINPUT14), .A3(G107), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G128), .B(G143), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n330), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n431), .A2(KEYINPUT14), .A3(G107), .A4(new_n436), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n290), .A2(G128), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G134), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n443), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n442), .A2(new_n447), .A3(G134), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n438), .A3(new_n450), .A4(new_n439), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n268), .A2(new_n259), .A3(new_n188), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT98), .A3(new_n252), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT98), .B1(new_n457), .B2(new_n252), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n458), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n428), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT91), .Z(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n429), .A2(G119), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT68), .B(G116), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n472), .B2(new_n208), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT2), .B(G113), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n283), .C1(new_n300), .C2(new_n301), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n473), .A2(new_n474), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n471), .A2(KEYINPUT5), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n470), .B1(new_n435), .B2(G119), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(KEYINPUT5), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n477), .B1(new_n480), .B2(G113), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n327), .ZN(new_n482));
  AOI211_X1 g296(.A(KEYINPUT6), .B(new_n469), .C1(new_n476), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n322), .A2(new_n194), .A3(new_n308), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n295), .A2(G125), .A3(new_n296), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(G224), .B2(new_n188), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n188), .A2(G224), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n484), .B2(new_n485), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n476), .A2(new_n482), .A3(new_n469), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n476), .A2(new_n482), .A3(new_n493), .A4(new_n469), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n469), .B1(new_n476), .B2(new_n482), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n483), .B(new_n490), .C1(new_n495), .C2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n481), .B1(new_n500), .B2(KEYINPUT90), .ZN(new_n501));
  INV_X1    g315(.A(new_n478), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(G113), .C1(new_n503), .C2(new_n473), .ZN(new_n504));
  INV_X1    g318(.A(new_n477), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n327), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n469), .B(KEYINPUT8), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n501), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n488), .A2(KEYINPUT7), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n486), .B(new_n512), .Z(new_n513));
  NAND3_X1  g327(.A1(new_n495), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n252), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n468), .B1(new_n499), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n495), .A2(new_n498), .ZN(new_n517));
  INV_X1    g331(.A(new_n483), .ZN(new_n518));
  INV_X1    g332(.A(new_n490), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n510), .B1(new_n492), .B2(new_n494), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n521), .B2(new_n513), .ZN(new_n522));
  INV_X1    g336(.A(new_n468), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G214), .B1(G237), .B2(G902), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT88), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n188), .A2(G952), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(G234), .B2(G237), .ZN(new_n530));
  OAI211_X1 g344(.A(G902), .B(G953), .C1(new_n260), .C2(new_n388), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT99), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT21), .B(G898), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n466), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n330), .A2(G137), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n332), .A2(G134), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n339), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n342), .A2(new_n297), .B1(new_n359), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n475), .B1(new_n541), .B2(KEYINPUT70), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n359), .A2(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n297), .A2(new_n341), .A3(new_n340), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT70), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT28), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT71), .ZN(new_n548));
  INV_X1    g362(.A(new_n475), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n297), .A2(new_n341), .A3(new_n340), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n539), .B1(new_n322), .B2(new_n308), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n475), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n547), .A2(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n388), .A2(new_n188), .A3(G210), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n298), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n558), .B(new_n559), .Z(new_n560));
  AOI211_X1 g374(.A(new_n548), .B(new_n555), .C1(new_n550), .C2(new_n553), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n556), .A2(KEYINPUT29), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n564));
  INV_X1    g378(.A(new_n560), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n543), .A2(KEYINPUT70), .A3(new_n544), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n549), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n555), .B1(new_n567), .B2(new_n545), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n551), .A2(new_n475), .A3(new_n552), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT66), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n539), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n540), .A2(KEYINPUT66), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n359), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n549), .B1(new_n573), .B2(new_n544), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT28), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n565), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT30), .B1(new_n551), .B2(new_n552), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n578), .A3(new_n544), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n549), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n580), .A2(new_n569), .A3(new_n560), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n564), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n563), .A2(new_n252), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT72), .A3(G472), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT72), .B1(new_n583), .B2(G472), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT32), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n573), .A2(new_n578), .A3(new_n544), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n578), .B1(new_n543), .B2(new_n544), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n475), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT69), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT31), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n590), .A2(new_n550), .A3(new_n560), .A4(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(KEYINPUT31), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n580), .A2(new_n569), .ZN(new_n596));
  INV_X1    g410(.A(new_n594), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(new_n560), .A3(new_n592), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n568), .A2(new_n575), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n565), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G472), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n587), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n595), .A2(new_n598), .B1(new_n600), .B2(new_n565), .ZN(new_n605));
  NOR4_X1   g419(.A1(new_n605), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n585), .A2(new_n586), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n387), .A2(new_n535), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n599), .A2(new_n601), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n252), .ZN(new_n611));
  NAND2_X1  g425(.A1(KEYINPUT100), .A2(G472), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n387), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n457), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n454), .A2(KEYINPUT33), .A3(new_n456), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n459), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n457), .A2(new_n459), .A3(new_n252), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n459), .A2(new_n252), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n427), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n516), .A2(new_n626), .A3(new_n524), .ZN(new_n627));
  INV_X1    g441(.A(new_n526), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n523), .B1(new_n520), .B2(new_n522), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(KEYINPUT102), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n627), .A2(new_n630), .A3(KEYINPUT103), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n627), .B2(new_n630), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n631), .A2(new_n632), .A3(new_n534), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n615), .A2(new_n625), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(G6));
  XOR2_X1   g451(.A(new_n426), .B(KEYINPUT105), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n464), .A2(new_n421), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n615), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT106), .Z(new_n645));
  OR3_X1    g459(.A1(new_n249), .A2(new_n250), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n645), .B1(new_n249), .B2(new_n250), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n646), .A2(new_n647), .A3(new_n265), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n258), .B2(new_n262), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n386), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n535), .A2(new_n650), .A3(new_n613), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  OAI21_X1  g467(.A(KEYINPUT32), .B1(new_n611), .B2(G472), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n602), .A2(new_n587), .A3(new_n603), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n582), .A2(new_n252), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n555), .B1(new_n550), .B2(new_n553), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n568), .B2(KEYINPUT71), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n658), .A2(new_n561), .A3(new_n564), .A4(new_n565), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT72), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n654), .A2(new_n655), .B1(new_n662), .B2(new_n584), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n520), .A2(new_n523), .A3(new_n522), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n629), .A3(KEYINPUT102), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n526), .B1(new_n516), .B2(new_n626), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n627), .A2(new_n630), .A3(KEYINPUT103), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n530), .B1(new_n532), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n638), .A2(new_n639), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n671), .A2(KEYINPUT107), .A3(new_n650), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n631), .A2(new_n632), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n650), .A3(new_n607), .A4(new_n674), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  INV_X1    g495(.A(new_n386), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n673), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  INV_X1    g499(.A(new_n649), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n654), .A2(new_n655), .ZN(new_n687));
  INV_X1    g501(.A(new_n554), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n252), .B1(new_n688), .B2(new_n560), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n596), .A2(new_n565), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n686), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n685), .A2(new_n526), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n428), .A2(new_n465), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n525), .B(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n694), .B(new_n696), .C1(new_n684), .C2(KEYINPUT40), .ZN(new_n697));
  OR3_X1    g511(.A1(new_n693), .A2(KEYINPUT109), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT109), .B1(new_n693), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n290), .ZN(G45));
  INV_X1    g515(.A(new_n673), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n427), .A2(new_n623), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n676), .A2(new_n650), .A3(new_n607), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NAND2_X1  g520(.A1(new_n662), .A2(new_n584), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n267), .B1(new_n687), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n273), .A2(KEYINPUT110), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n380), .A2(new_n381), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n709), .B1(new_n710), .B2(G902), .ZN(new_n711));
  OAI221_X1 g525(.A(new_n252), .B1(KEYINPUT110), .B2(new_n273), .C1(new_n380), .C2(new_n381), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n272), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n633), .A3(new_n625), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NOR3_X1   g531(.A1(new_n631), .A2(new_n632), .A3(new_n713), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n258), .A2(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n640), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n534), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n607), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NOR2_X1   g537(.A1(new_n649), .A2(new_n466), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n718), .A2(new_n721), .A3(new_n607), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NOR3_X1   g540(.A1(new_n713), .A2(new_n428), .A3(new_n465), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n603), .A2(new_n252), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n556), .A2(new_n562), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n565), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n730), .B2(new_n599), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n611), .B2(G472), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(new_n719), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n732), .B2(new_n719), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n633), .B(new_n727), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  AOI22_X1  g551(.A1(new_n729), .A2(new_n565), .B1(new_n595), .B2(new_n598), .ZN(new_n738));
  OAI22_X1  g552(.A1(new_n602), .A2(new_n603), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n649), .A2(new_n739), .A3(new_n703), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n676), .A3(new_n714), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  OAI211_X1 g556(.A(new_n382), .B(new_n384), .C1(new_n273), .C2(new_n366), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(new_n272), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n525), .A2(new_n628), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n708), .A2(new_n704), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n708), .A2(new_n746), .A3(KEYINPUT42), .A4(new_n704), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  AND3_X1   g566(.A1(new_n708), .A2(new_n746), .A3(new_n674), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n330), .ZN(G36));
  INV_X1    g568(.A(new_n745), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n428), .A2(new_n756), .A3(new_n623), .ZN(new_n757));
  OR3_X1    g571(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n758), .B2(new_n427), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OR3_X1    g574(.A1(new_n760), .A2(new_n613), .A3(new_n649), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n761), .A2(KEYINPUT113), .A3(new_n762), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n755), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n761), .A2(new_n762), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n367), .A2(new_n769), .A3(new_n378), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n384), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n382), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT112), .B1(new_n773), .B2(new_n382), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n772), .B2(new_n384), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n271), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n767), .A2(new_n683), .A3(new_n768), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n777), .B2(new_n271), .ZN(new_n782));
  INV_X1    g596(.A(new_n775), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n382), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT47), .B(new_n272), .C1(new_n785), .C2(new_n776), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n607), .A2(new_n719), .A3(new_n703), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n745), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND2_X1  g604(.A1(new_n711), .A2(new_n712), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT49), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT114), .Z(new_n793));
  AOI211_X1 g607(.A(new_n271), .B(new_n793), .C1(KEYINPUT49), .C2(new_n791), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n687), .A2(new_n719), .A3(new_n691), .ZN(new_n795));
  INV_X1    g609(.A(new_n527), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n795), .A2(new_n796), .A3(new_n696), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n428), .A3(new_n623), .A4(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n705), .A2(new_n741), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n670), .A2(new_n428), .A3(new_n465), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n702), .A3(new_n692), .A4(new_n744), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n677), .A2(new_n678), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n677), .A2(new_n678), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n799), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n705), .A2(new_n741), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n675), .B2(new_n679), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n801), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n805), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(new_n805), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n428), .A2(new_n464), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n528), .B1(new_n815), .B2(new_n624), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n387), .A2(new_n816), .A3(new_n721), .A4(new_n613), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n736), .A2(new_n725), .A3(new_n608), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n715), .A2(new_n722), .A3(new_n651), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n753), .B1(new_n749), .B2(new_n750), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n746), .A2(new_n740), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n638), .A2(new_n673), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n650), .A2(new_n421), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n465), .A3(new_n607), .A4(new_n745), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT53), .A4(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n809), .A2(new_n680), .A3(new_n799), .A4(new_n801), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n809), .B1(new_n808), .B2(new_n801), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n805), .A2(new_n806), .A3(new_n810), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n805), .A2(new_n810), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(new_n826), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(KEYINPUT116), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n837), .A3(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(new_n530), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n714), .A2(new_n745), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n795), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n625), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n831), .A2(new_n834), .A3(new_n827), .A4(new_n832), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT53), .B1(new_n835), .B2(new_n826), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT54), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n757), .A2(new_n530), .A3(new_n759), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT117), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n734), .A2(new_n735), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n718), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n849), .A2(new_n714), .A3(new_n745), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n686), .A3(new_n732), .ZN(new_n854));
  NAND2_X1  g668(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n855));
  NOR2_X1   g669(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n713), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n696), .A2(new_n526), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n851), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n849), .A2(new_n850), .A3(new_n858), .ZN(new_n860));
  OAI211_X1 g674(.A(KEYINPUT118), .B(KEYINPUT50), .C1(new_n860), .C2(new_n713), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n841), .A2(new_n428), .A3(new_n758), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n854), .A2(new_n859), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n791), .A2(new_n272), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n782), .A2(new_n786), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n851), .A2(new_n745), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT51), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n529), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n782), .A2(new_n786), .A3(new_n872), .A4(new_n865), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n867), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT51), .A3(new_n863), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n852), .B(new_n870), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n853), .A2(new_n708), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT48), .Z(new_n881));
  NOR3_X1   g695(.A1(new_n847), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(G952), .A2(G953), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n798), .B1(new_n882), .B2(new_n883), .ZN(G75));
  NAND4_X1  g698(.A1(new_n843), .A2(G902), .A3(new_n468), .A4(new_n844), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n517), .A2(new_n518), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n490), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n520), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT55), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n188), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n891), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n885), .A2(new_n886), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n892), .A2(new_n899), .A3(new_n894), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(new_n383), .B(KEYINPUT57), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n845), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n710), .B(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n843), .A2(new_n844), .ZN(new_n907));
  OR3_X1    g721(.A1(new_n907), .A2(new_n252), .A3(new_n772), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n893), .B1(new_n906), .B2(new_n908), .ZN(G54));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n252), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n410), .A2(new_n415), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n893), .ZN(G60));
  AND2_X1   g730(.A1(new_n617), .A2(new_n618), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n622), .B(KEYINPUT59), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n919), .C1(new_n903), .C2(new_n845), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n838), .B2(new_n846), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n920), .B(new_n894), .C1(new_n921), .C2(new_n917), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(G217), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n252), .ZN(new_n926));
  NAND3_X1  g740(.A1(KEYINPUT60), .A2(G217), .A3(G902), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n646), .A2(new_n647), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT123), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n843), .A2(new_n844), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n907), .B1(new_n926), .B2(new_n927), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n894), .B(new_n931), .C1(new_n932), .C2(new_n264), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n894), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT61), .B1(new_n934), .B2(KEYINPUT124), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G66));
  INV_X1    g750(.A(G224), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n533), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n820), .B2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n888), .B1(G898), .B2(new_n188), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  NAND2_X1  g755(.A1(new_n577), .A2(new_n579), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n412), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n779), .A2(new_n789), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n821), .A3(new_n808), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n683), .A2(new_n778), .A3(new_n708), .A4(new_n800), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n188), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n672), .A2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n951));
  INV_X1    g765(.A(new_n943), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n698), .A2(new_n699), .A3(new_n808), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n684), .B1(new_n624), .B2(new_n815), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n708), .A3(new_n745), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n944), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n952), .B1(new_n958), .B2(new_n188), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n950), .A2(new_n951), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n951), .B1(new_n950), .B2(new_n959), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G72));
  XNOR2_X1  g776(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n603), .A2(new_n252), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n945), .A2(new_n946), .ZN(new_n966));
  INV_X1    g780(.A(new_n820), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n581), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n958), .B2(new_n967), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n893), .B1(new_n970), .B2(new_n690), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n690), .A2(new_n581), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n828), .A2(new_n837), .A3(new_n965), .A4(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(G57));
endmodule


