//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT11), .A2(G134), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT65), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT65), .A2(G137), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n195), .B(new_n189), .C1(new_n191), .C2(new_n192), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT67), .B(G131), .Z(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT11), .A2(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n188), .B1(new_n199), .B2(G137), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n196), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G134), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n203), .B(KEYINPUT69), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n191), .A2(new_n192), .A3(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(G131), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT70), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT1), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT71), .B(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n220), .A2(new_n211), .A3(new_n216), .A4(G128), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n201), .B(new_n206), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT64), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n217), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(KEYINPUT0), .A3(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n225), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n202), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n188), .B1(new_n236), .B2(new_n190), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n200), .B1(new_n237), .B2(new_n195), .ZN(new_n238));
  INV_X1    g052(.A(new_n196), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n240), .B2(new_n201), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n222), .B1(new_n241), .B2(KEYINPUT68), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  AOI211_X1 g057(.A(new_n243), .B(new_n234), .C1(new_n240), .C2(new_n201), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n187), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT72), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT2), .B(G113), .Z(new_n247));
  XNOR2_X1  g061(.A(G116), .B(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G116), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(G116), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n255), .A3(KEYINPUT73), .ZN(new_n256));
  OR3_X1    g070(.A1(new_n247), .A2(KEYINPUT73), .A3(new_n248), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(new_n187), .C1(new_n242), .C2(new_n244), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n240), .A2(new_n201), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n225), .A2(new_n232), .A3(new_n233), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n264), .A2(new_n222), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT30), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n246), .A2(new_n259), .A3(new_n261), .A4(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n264), .A2(new_n258), .A3(new_n222), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G237), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G210), .ZN(new_n272));
  INV_X1    g086(.A(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND3_X1  g090(.A1(new_n267), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT31), .ZN(new_n278));
  INV_X1    g092(.A(new_n276), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n259), .B1(new_n242), .B2(new_n244), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n268), .B1(new_n281), .B2(KEYINPUT74), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n283), .B(new_n259), .C1(new_n242), .C2(new_n244), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n268), .A2(KEYINPUT28), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n279), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n267), .A2(new_n288), .A3(new_n269), .A4(new_n276), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n278), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n285), .A2(new_n286), .A3(new_n279), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n276), .B1(new_n267), .B2(new_n269), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(KEYINPUT29), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n286), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n265), .A2(new_n258), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n268), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n298), .B(new_n299), .C1(new_n301), .C2(new_n280), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n303), .B2(new_n302), .ZN(new_n305));
  OAI21_X1  g119(.A(G472), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(G113), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(new_n248), .B2(new_n247), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G107), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G104), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n273), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(G104), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n316), .B2(G107), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(KEYINPUT3), .A3(G104), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n320), .B1(new_n325), .B2(new_n273), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n315), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n325), .B2(new_n273), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n318), .A2(KEYINPUT3), .A3(G104), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT3), .B1(new_n318), .B2(G104), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n317), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G101), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n331), .A3(G101), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n257), .A3(new_n256), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G122), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n330), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n234), .A2(G125), .ZN(new_n342));
  INV_X1    g156(.A(G125), .ZN(new_n343));
  INV_X1    g157(.A(new_n221), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n218), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT87), .B(G224), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n271), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT7), .A4(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n340), .B(KEYINPUT8), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n325), .A2(new_n273), .ZN(new_n351));
  INV_X1    g165(.A(new_n320), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n315), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n313), .A2(new_n314), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n249), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n326), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n347), .B1(new_n342), .B2(new_n345), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT7), .B1(new_n342), .B2(new_n345), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n349), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n340), .ZN(new_n363));
  INV_X1    g177(.A(new_n339), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(KEYINPUT85), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n326), .A2(new_n327), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n356), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n342), .A2(new_n345), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(new_n347), .Z(new_n371));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(new_n363), .C1(new_n364), .C2(new_n367), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G210), .B1(G237), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n362), .A2(new_n374), .A3(new_n376), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n310), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(KEYINPUT9), .B(G234), .Z(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G221), .B1(new_n382), .B2(G902), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n263), .A2(new_n337), .A3(new_n338), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT82), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n263), .A2(new_n337), .A3(new_n386), .A4(new_n338), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n208), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n211), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(G128), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n221), .B1(new_n393), .B2(new_n217), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n389), .B1(new_n394), .B2(new_n353), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT84), .B(new_n389), .C1(new_n394), .C2(new_n353), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n262), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n365), .A2(new_n366), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n389), .B1(new_n218), .B2(new_n344), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n388), .A2(new_n399), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n271), .A2(G227), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n405), .B(new_n406), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(KEYINPUT86), .A3(new_n407), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n219), .A2(new_n221), .A3(new_n326), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n394), .A2(new_n353), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n262), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT12), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT12), .B(new_n262), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n410), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n388), .A2(new_n399), .A3(new_n403), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n262), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n404), .ZN(new_n422));
  INV_X1    g236(.A(new_n407), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI211_X1 g238(.A(G469), .B(G902), .C1(new_n419), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n404), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n423), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n404), .A3(new_n407), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G902), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n380), .B(new_n383), .C1(new_n425), .C2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n381), .A2(G217), .A3(new_n271), .ZN(new_n434));
  INV_X1    g248(.A(G122), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n318), .B1(new_n436), .B2(KEYINPUT14), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n226), .A2(KEYINPUT71), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G143), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n226), .A2(G143), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n441), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n207), .B1(new_n442), .B2(new_n444), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(KEYINPUT95), .A3(new_n447), .ZN(new_n451));
  OAI21_X1  g265(.A(G134), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT95), .B1(new_n450), .B2(new_n447), .ZN(new_n453));
  INV_X1    g267(.A(G134), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n441), .B(new_n448), .C1(new_n214), .C2(new_n207), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n440), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n448), .B(new_n458), .C1(new_n214), .C2(new_n207), .ZN(new_n459));
  AND2_X1   g273(.A1(KEYINPUT94), .A2(KEYINPUT13), .ZN(new_n460));
  NOR2_X1   g274(.A1(KEYINPUT94), .A2(KEYINPUT13), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n454), .B1(new_n462), .B2(new_n447), .ZN(new_n463));
  XOR2_X1   g277(.A(G116), .B(G122), .Z(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G107), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n438), .A2(new_n318), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n459), .A2(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n456), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n434), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n439), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n434), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n468), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n474), .A2(KEYINPUT96), .A3(new_n468), .A4(new_n475), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G478), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n479), .A2(KEYINPUT97), .A3(new_n431), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n431), .A3(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT97), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT98), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n483), .B(new_n490), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G125), .B(G140), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT16), .ZN(new_n494));
  OR3_X1    g308(.A1(new_n343), .A2(KEYINPUT16), .A3(G140), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n210), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(G146), .A3(new_n495), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT91), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G214), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n504), .A2(G237), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(G143), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(G143), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n197), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n198), .B(new_n507), .C1(new_n505), .C2(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT92), .B1(new_n512), .B2(KEYINPUT17), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(KEYINPUT17), .A3(new_n197), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n510), .A2(new_n515), .A3(new_n516), .A4(new_n511), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n503), .A2(new_n513), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n493), .A2(new_n210), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT78), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n210), .B2(new_n493), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n509), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT90), .B(G104), .Z(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT93), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n518), .A2(KEYINPUT93), .A3(new_n529), .A4(new_n524), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n431), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G475), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(G952), .A3(new_n271), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT21), .B(G898), .Z(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(G902), .A3(G953), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n529), .B1(new_n518), .B2(new_n524), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n493), .B(KEYINPUT19), .Z(new_n546));
  OAI21_X1  g360(.A(new_n498), .B1(new_n546), .B2(G146), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT89), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n498), .C1(new_n546), .C2(G146), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n512), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n528), .B1(new_n521), .B2(new_n523), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G475), .A2(G902), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n544), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  NOR4_X1   g371(.A1(new_n545), .A2(new_n553), .A3(KEYINPUT20), .A4(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n534), .B(new_n543), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n492), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n433), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(KEYINPUT24), .A2(G110), .ZN(new_n563));
  NAND2_X1  g377(.A1(KEYINPUT24), .A2(G110), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT76), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n226), .A2(G119), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n214), .B2(new_n251), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT77), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT23), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n226), .A3(G119), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n572), .B2(new_n575), .ZN(new_n577));
  INV_X1    g391(.A(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n569), .A2(new_n580), .A3(new_n572), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n520), .A2(new_n498), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n577), .A2(new_n578), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n569), .A2(new_n572), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n499), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT22), .B(G137), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n271), .A2(G221), .A3(G234), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n584), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n499), .A2(new_n586), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n585), .A2(new_n593), .B1(new_n582), .B2(new_n583), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n590), .B(KEYINPUT79), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n592), .B(new_n431), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n584), .A2(new_n587), .ZN(new_n599));
  INV_X1    g413(.A(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n601), .A2(new_n431), .A3(new_n592), .A4(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G217), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(G234), .B2(new_n431), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT81), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT81), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n598), .A2(new_n609), .A3(new_n604), .A4(new_n606), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n601), .A2(new_n592), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n606), .A2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n308), .A2(new_n562), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT99), .B(G101), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G3));
  NAND2_X1  g432(.A1(new_n290), .A2(new_n431), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n620), .A2(new_n292), .ZN(new_n621));
  INV_X1    g435(.A(new_n383), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n419), .A2(new_n424), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n426), .A3(new_n431), .ZN(new_n624));
  INV_X1    g438(.A(new_n432), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n615), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n380), .A2(new_n543), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n534), .B1(new_n556), .B2(new_n558), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n479), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n470), .A2(KEYINPUT33), .A3(new_n476), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(G478), .A3(new_n431), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n484), .A2(new_n480), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n633), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT100), .B1(new_n641), .B2(new_n630), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NOR3_X1   g460(.A1(new_n492), .A2(new_n630), .A3(new_n633), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n629), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n600), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n599), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n612), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n608), .A2(new_n610), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n620), .A2(new_n292), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n620), .A2(KEYINPUT101), .A3(new_n292), .A4(new_n654), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n562), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(new_n433), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n537), .B1(new_n541), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n492), .A2(new_n633), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n308), .A2(new_n663), .A3(new_n654), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT103), .B(G128), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G30));
  XNOR2_X1  g483(.A(new_n665), .B(KEYINPUT39), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n626), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT40), .Z(new_n673));
  AOI21_X1  g487(.A(new_n279), .B1(new_n267), .B2(new_n269), .ZN(new_n674));
  AOI21_X1  g488(.A(G902), .B1(new_n301), .B2(new_n279), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n294), .A2(new_n307), .A3(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n489), .A2(new_n491), .ZN(new_n679));
  INV_X1    g493(.A(new_n654), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n309), .A3(new_n633), .A4(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n378), .A2(new_n379), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT38), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n681), .B2(KEYINPUT104), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n673), .A2(new_n678), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NOR2_X1   g502(.A1(new_n641), .A2(new_n665), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n308), .A2(new_n663), .A3(new_n654), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AOI22_X1  g505(.A1(new_n408), .A2(new_n409), .B1(new_n417), .B2(new_n416), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n692), .A2(new_n411), .B1(new_n422), .B2(new_n423), .ZN(new_n693));
  OAI21_X1  g507(.A(G469), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n624), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n622), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n643), .A2(new_n308), .A3(new_n615), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n308), .A2(new_n615), .A3(new_n647), .A4(new_n696), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n561), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n426), .B1(new_n623), .B2(new_n431), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n425), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n380), .A4(new_n383), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n624), .A3(new_n380), .A4(new_n383), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT105), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND4_X1   g523(.A1(new_n702), .A2(new_n709), .A3(new_n308), .A4(new_n654), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n251), .ZN(G21));
  NOR2_X1   g525(.A1(new_n301), .A2(new_n280), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n279), .B1(new_n712), .B2(new_n286), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n278), .A2(new_n289), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n291), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n620), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n615), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n695), .A2(new_n622), .A3(new_n542), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n489), .A2(new_n380), .A3(new_n491), .A4(new_n633), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n435), .ZN(G24));
  AND4_X1   g539(.A1(new_n620), .A2(new_n654), .A3(new_n689), .A4(new_n715), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n709), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(new_n307), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT32), .B1(new_n290), .B2(new_n291), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n614), .B1(new_n731), .B2(new_n306), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n683), .A2(new_n310), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n626), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n689), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n308), .A2(new_n734), .A3(new_n615), .A4(new_n689), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  AND4_X1   g556(.A1(new_n308), .A2(new_n734), .A3(new_n615), .A4(new_n666), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n454), .ZN(G36));
  INV_X1    g558(.A(new_n633), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n639), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n621), .A2(new_n680), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n430), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n428), .A2(KEYINPUT45), .A3(new_n429), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(G469), .A2(G902), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT46), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n425), .B1(new_n766), .B2(KEYINPUT46), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n622), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n760), .A2(new_n671), .A3(new_n733), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n758), .A2(new_n759), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n202), .ZN(G39));
  NOR2_X1   g587(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n769), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n689), .A2(new_n733), .A3(new_n614), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n776), .A2(new_n779), .A3(new_n308), .A4(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(G140), .Z(G42));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n783));
  INV_X1    g597(.A(new_n717), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n536), .B1(new_n751), .B2(new_n752), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n684), .A2(new_n695), .A3(new_n309), .A4(new_n622), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI22_X1  g605(.A1(new_n776), .A2(new_n779), .B1(new_n383), .B2(new_n695), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n733), .A3(new_n787), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n696), .A2(new_n733), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n294), .A2(new_n307), .A3(new_n677), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n537), .A4(new_n615), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n633), .A3(new_n639), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n785), .A2(new_n795), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n785), .A2(new_n802), .A3(new_n795), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n716), .A2(new_n654), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(KEYINPUT116), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n799), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n783), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n808), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n798), .B1(new_n811), .B2(new_n806), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n791), .A4(new_n793), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n804), .A2(new_n732), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT48), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(G952), .B(new_n271), .C1(new_n797), .C2(new_n641), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n709), .B2(new_n787), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n814), .A2(new_n815), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n816), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n814), .A2(new_n815), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n810), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT118), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n743), .B1(new_n737), .B2(new_n740), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n745), .A2(new_n488), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n630), .B1(new_n828), .B2(new_n641), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n627), .A2(new_n292), .A3(new_n620), .A4(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n616), .B(new_n830), .C1(new_n717), .C2(new_n723), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n710), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n697), .A2(new_n659), .A3(new_n700), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n308), .A2(new_n654), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n633), .A2(new_n488), .A3(new_n665), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT112), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n734), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n835), .A2(new_n838), .B1(new_n726), .B2(new_n734), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n827), .A2(new_n832), .A3(new_n833), .A4(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n727), .A2(new_n667), .A3(new_n690), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n624), .A2(new_n625), .ZN(new_n843));
  INV_X1    g657(.A(new_n665), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n610), .A2(new_n608), .A3(new_n653), .A4(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n843), .A2(new_n845), .A3(new_n383), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n721), .B2(new_n722), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n842), .B1(new_n847), .B2(new_n796), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n626), .A2(new_n845), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n679), .A2(KEYINPUT106), .A3(new_n380), .A4(new_n633), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n719), .A2(new_n720), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(KEYINPUT113), .A3(new_n678), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n854), .A3(KEYINPUT52), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n847), .A2(new_n796), .A3(new_n842), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT113), .B1(new_n852), .B2(new_n678), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n727), .A2(new_n667), .A3(new_n690), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n841), .B2(new_n854), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n856), .A3(new_n855), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n840), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(KEYINPUT53), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n827), .A2(new_n832), .A3(new_n833), .A4(new_n839), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n855), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT54), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n869), .B2(new_n870), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n867), .B2(KEYINPUT53), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n826), .A2(new_n879), .B1(G952), .B2(G953), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n695), .A2(KEYINPUT49), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT111), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n695), .A2(KEYINPUT49), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n615), .A2(new_n309), .A3(new_n383), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n884), .A2(new_n684), .A3(new_n885), .A4(new_n746), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(KEYINPUT111), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n880), .B1(new_n678), .B2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n271), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n876), .A2(new_n431), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n369), .A2(new_n373), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n371), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n891), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n865), .B1(new_n856), .B2(new_n855), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n841), .C2(new_n854), .ZN(new_n899));
  OAI211_X1 g713(.A(KEYINPUT53), .B(new_n869), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n871), .A2(new_n872), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT119), .B1(new_n902), .B2(G902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n431), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n377), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n896), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n897), .B1(new_n908), .B2(new_n910), .ZN(G51));
  AOI21_X1  g725(.A(KEYINPUT120), .B1(new_n902), .B2(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n878), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n876), .A2(KEYINPUT120), .A3(new_n877), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n765), .B(KEYINPUT57), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n693), .B(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n906), .A2(new_n764), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n890), .B1(new_n918), .B2(new_n919), .ZN(G54));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n904), .B1(new_n876), .B2(new_n431), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n902), .A2(KEYINPUT119), .A3(G902), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n891), .B1(new_n925), .B2(new_n554), .ZN(new_n926));
  INV_X1    g740(.A(new_n554), .ZN(new_n927));
  AOI211_X1 g741(.A(new_n927), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n921), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n906), .B2(new_n922), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n554), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT122), .A4(new_n891), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(G60));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n874), .B2(new_n878), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n635), .A2(new_n636), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n891), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n913), .A2(new_n914), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n937), .A2(new_n935), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT124), .ZN(new_n944));
  XOR2_X1   g758(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n876), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n652), .B(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n891), .C1(new_n611), .C2(new_n947), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G66));
  AOI21_X1  g766(.A(new_n271), .B1(new_n538), .B2(new_n346), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n832), .A2(new_n833), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n271), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n894), .B1(G898), .B2(new_n271), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT126), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  NAND3_X1  g772(.A1(new_n246), .A2(new_n261), .A3(new_n266), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT127), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n546), .ZN(new_n961));
  OAI211_X1 g775(.A(G900), .B(G953), .C1(new_n961), .C2(G227), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(G227), .B2(new_n961), .ZN(new_n963));
  INV_X1    g777(.A(new_n732), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n769), .B(new_n671), .C1(new_n721), .C2(new_n722), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n827), .B(new_n841), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n772), .A2(new_n966), .A3(new_n781), .ZN(new_n967));
  INV_X1    g781(.A(new_n961), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(G953), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n772), .A2(new_n781), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n687), .A2(new_n841), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n828), .A2(new_n641), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n733), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n964), .A2(new_n672), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n971), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n968), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n963), .B1(new_n970), .B2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n977), .B2(new_n954), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n674), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n267), .A2(new_n269), .A3(new_n279), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n967), .A2(new_n954), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n981), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n868), .A2(new_n873), .ZN(new_n987));
  INV_X1    g801(.A(new_n277), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n988), .B2(new_n296), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n983), .A2(new_n986), .A3(new_n890), .A4(new_n990), .ZN(G57));
endmodule


