//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n211), .B1(new_n212), .B2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n214), .A2(KEYINPUT66), .A3(G1), .A4(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n219), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G68), .B2(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  INV_X1    g0029(.A(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G77), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n201), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n212), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NAND2_X1  g0037(.A1(G1), .A2(G13), .ZN(new_n238));
  INV_X1    g0038(.A(G20), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n206), .A2(new_n229), .ZN(new_n241));
  AOI211_X1 g0041(.A(new_n218), .B(new_n237), .C1(new_n240), .C2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n226), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n229), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n201), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  OR2_X1    g0057(.A1(KEYINPUT68), .A2(G58), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT68), .A2(G58), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n258), .B(KEYINPUT8), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n259), .A2(new_n201), .A3(KEYINPUT8), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n239), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n265), .B1(G150), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n208), .A2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n270), .A2(KEYINPUT67), .A3(new_n238), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT67), .B1(new_n270), .B2(new_n238), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n214), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n269), .A2(new_n273), .B1(new_n229), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n270), .A2(new_n238), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n270), .A2(KEYINPUT67), .A3(new_n238), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G50), .A3(new_n275), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OR2_X1    g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G222), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G223), .A2(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n295), .B(new_n298), .C1(G77), .C2(new_n291), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n274), .B(G274), .C1(G41), .C2(G45), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n299), .B(new_n300), .C1(new_n230), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT72), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G200), .B2(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n288), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT10), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(G179), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n303), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n284), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n230), .A2(new_n292), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n291), .B(new_n316), .C1(G232), .C2(new_n292), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n297), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n297), .A2(G238), .A3(new_n301), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n300), .B(KEYINPUT73), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n322), .ZN(new_n324));
  NOR4_X1   g0124(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT13), .A4(new_n320), .ZN(new_n325));
  OAI21_X1  g0125(.A(G169), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n323), .A2(new_n325), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G179), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(G169), .C1(new_n323), .C2(new_n325), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n231), .B2(new_n264), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n273), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n336));
  XOR2_X1   g0136(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g0137(.A(new_n275), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n278), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G68), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n276), .A2(new_n202), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n341), .A2(KEYINPUT12), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(KEYINPUT12), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n337), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n332), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G238), .A2(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n291), .B(new_n346), .C1(new_n234), .C2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n298), .C1(G107), .C2(new_n291), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n300), .C1(new_n232), .C2(new_n302), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT70), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT70), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n349), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n311), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n264), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n278), .B1(new_n231), .B2(new_n276), .ZN(new_n361));
  INV_X1    g0161(.A(new_n339), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n231), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n352), .A2(new_n355), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n345), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT77), .ZN(new_n368));
  INV_X1    g0168(.A(new_n300), .ZN(new_n369));
  OR2_X1    g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n230), .A2(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(new_n290), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n376), .B2(new_n298), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n297), .A2(G232), .A3(new_n301), .ZN(new_n378));
  AOI21_X1  g0178(.A(G200), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n297), .B1(new_n374), .B2(new_n375), .ZN(new_n380));
  INV_X1    g0180(.A(new_n378), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n380), .A2(new_n381), .A3(G190), .A4(new_n369), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n368), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(new_n304), .A3(new_n378), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n380), .A2(new_n381), .A3(new_n369), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(KEYINPUT77), .C1(G200), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(KEYINPUT68), .A2(G58), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT68), .A2(G58), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n206), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT75), .B(G68), .C1(new_n388), .C2(new_n389), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G20), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n372), .A2(new_n373), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n397), .B2(new_n239), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NOR4_X1   g0199(.A1(new_n372), .A2(new_n373), .A3(new_n399), .A4(G20), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n266), .A2(G159), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n401), .A4(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n278), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n338), .A2(G13), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n263), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n263), .A2(new_n275), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT76), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n410), .B(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(new_n282), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n387), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n387), .A2(new_n407), .A3(KEYINPUT17), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n407), .A2(new_n413), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n385), .A2(new_n311), .ZN(new_n419));
  NOR4_X1   g0219(.A1(new_n380), .A2(new_n381), .A3(new_n351), .A4(new_n369), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n424), .B(new_n421), .C1(new_n407), .C2(new_n413), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n416), .B(new_n417), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n367), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n344), .B1(G190), .B2(new_n328), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n328), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n364), .B(new_n361), .C1(new_n350), .C2(new_n429), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n354), .A2(new_n304), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n314), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT6), .ZN(new_n437));
  AND2_X1   g0237(.A1(G97), .A2(G107), .ZN(new_n438));
  NOR2_X1   g0238(.A1(G97), .A2(G107), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n225), .A2(KEYINPUT6), .A3(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G20), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n266), .A2(G77), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n399), .B1(new_n291), .B2(G20), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n239), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n225), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n278), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n276), .A2(new_n221), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT78), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n274), .A2(G33), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n408), .B(new_n453), .C1(new_n271), .C2(new_n272), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n449), .B(new_n452), .C1(new_n456), .C2(new_n221), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT85), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G274), .A3(new_n297), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n274), .B(G45), .C1(new_n458), .C2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT83), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n461), .A2(G41), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT83), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT84), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT84), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n469), .A2(KEYINPUT83), .A3(new_n470), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n464), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n463), .A2(new_n473), .A3(new_n475), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n478), .A2(new_n297), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(G257), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G244), .B(new_n292), .C1(new_n372), .C2(new_n373), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT81), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n484), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n485), .B(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n220), .B1(new_n289), .B2(new_n290), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(G1698), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(KEYINPUT82), .A3(new_n483), .A4(new_n484), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n495), .A3(new_n298), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n480), .A2(new_n496), .A3(G179), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n311), .B1(new_n480), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n457), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n480), .A2(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G200), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n282), .A2(new_n455), .A3(new_n453), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n454), .A2(KEYINPUT79), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n221), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n270), .A2(new_n238), .ZN(new_n506));
  OAI21_X1  g0306(.A(G107), .B1(new_n398), .B2(new_n400), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n442), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT80), .B1(new_n510), .B2(new_n452), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  NOR4_X1   g0312(.A1(new_n505), .A2(new_n509), .A3(new_n512), .A4(new_n451), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n502), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n480), .A2(new_n496), .A3(G190), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n480), .A2(new_n496), .A3(KEYINPUT86), .A4(G190), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n500), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n463), .A2(G274), .A3(new_n297), .ZN(new_n523));
  INV_X1    g0323(.A(new_n476), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n291), .A2(G250), .A3(new_n292), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n291), .A2(G257), .A3(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(G33), .ZN(new_n529));
  INV_X1    g0329(.A(G294), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n298), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n478), .A2(G264), .A3(new_n297), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT92), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n478), .A2(KEYINPUT92), .A3(G264), .A4(new_n297), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(new_n526), .A3(new_n532), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n535), .B1(new_n540), .B2(new_n351), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n239), .B(G87), .C1(new_n372), .C2(new_n373), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n291), .A2(new_n544), .A3(new_n239), .A4(G87), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n543), .A2(new_n545), .B1(G116), .B2(new_n265), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n239), .A2(G107), .B1(KEYINPUT91), .B2(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g0347(.A1(KEYINPUT91), .A2(KEYINPUT23), .ZN(new_n548));
  XOR2_X1   g0348(.A(new_n547), .B(new_n548), .Z(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(KEYINPUT24), .A3(new_n549), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n278), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n276), .A2(new_n225), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n555), .B(KEYINPUT25), .Z(new_n556));
  NAND2_X1  g0356(.A1(new_n503), .A2(new_n504), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n541), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n540), .A2(new_n429), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n304), .A2(new_n526), .A3(new_n532), .A4(new_n533), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT93), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT93), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n562), .B1(new_n540), .B2(new_n429), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(new_n559), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n560), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n478), .A2(G270), .A3(new_n297), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n477), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(new_n292), .C1(new_n372), .C2(new_n373), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT89), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n291), .A2(KEYINPUT89), .A3(G257), .A4(new_n292), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n397), .A2(G303), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n291), .A2(G264), .A3(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT90), .A3(new_n298), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT90), .B1(new_n580), .B2(new_n298), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n573), .B(G190), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G116), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n276), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n408), .A2(G116), .A3(new_n506), .A4(new_n453), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n506), .B1(G20), .B2(new_n585), .ZN(new_n588));
  AOI21_X1  g0388(.A(G20), .B1(new_n529), .B2(G97), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n486), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n588), .A2(new_n590), .A3(KEYINPUT20), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n586), .B(new_n587), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n526), .A2(new_n571), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n580), .A2(new_n298), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n598), .B2(new_n581), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n584), .B(new_n594), .C1(new_n599), .C2(new_n429), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n593), .A2(G169), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(G179), .A3(new_n593), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n605), .A2(KEYINPUT21), .A3(G169), .A4(new_n593), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n600), .A2(new_n603), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n291), .B1(G244), .B2(new_n292), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G238), .A2(G1698), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(new_n529), .B2(new_n585), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n298), .ZN(new_n611));
  INV_X1    g0411(.A(G274), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n469), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n297), .C1(G250), .C2(new_n469), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(new_n429), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n439), .A2(new_n219), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n318), .A2(new_n239), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n264), .A2(KEYINPUT19), .A3(new_n221), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n291), .A2(new_n239), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(new_n202), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT88), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  OAI221_X1 g0425(.A(new_n625), .B1(new_n622), .B2(new_n202), .C1(new_n620), .C2(new_n621), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n626), .A3(new_n278), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n276), .A2(new_n359), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n615), .A2(G190), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n557), .A2(G87), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n616), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n351), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n456), .A2(new_n359), .ZN(new_n635));
  OAI221_X1 g0435(.A(new_n634), .B1(G169), .B2(new_n615), .C1(new_n629), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n607), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n457), .A2(new_n512), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n510), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n502), .A3(new_n517), .A4(new_n518), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(KEYINPUT87), .A3(new_n500), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n522), .A2(new_n570), .A3(new_n638), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n436), .A2(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n367), .A2(new_n430), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n416), .A2(new_n417), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n646), .A2(new_n647), .B1(new_n423), .B2(new_n425), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n309), .A2(new_n648), .B1(new_n284), .B2(new_n312), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n614), .B(KEYINPUT94), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n611), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n311), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n634), .B(new_n653), .C1(new_n629), .C2(new_n635), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n566), .A2(new_n569), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(G200), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n630), .A2(new_n631), .A3(new_n632), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n603), .A2(new_n606), .A3(new_n604), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n642), .B(new_n500), .C1(new_n661), .C2(new_n560), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n654), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n639), .B(new_n640), .C1(new_n498), .C2(new_n499), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n658), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT95), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n637), .ZN(new_n670));
  INV_X1    g0470(.A(new_n500), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(KEYINPUT26), .A3(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT95), .B(new_n665), .C1(new_n658), .C2(new_n666), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n650), .B1(new_n435), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT96), .Z(G369));
  NOR2_X1   g0477(.A1(new_n214), .A2(G20), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .A3(G1), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT27), .B1(new_n679), .B2(G1), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n570), .B1(new_n565), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n661), .A2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n560), .A2(new_n684), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n594), .A2(new_n685), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n661), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n607), .B2(new_n691), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n570), .A2(new_n687), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n560), .A2(new_n685), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n216), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n439), .A2(new_n219), .A3(new_n585), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n274), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n241), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  NOR3_X1   g0505(.A1(new_n637), .A2(KEYINPUT26), .A3(new_n500), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n658), .A2(new_n666), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(KEYINPUT26), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(new_n654), .C1(new_n660), .C2(new_n662), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n685), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n570), .A2(new_n638), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n522), .A3(new_n643), .A4(new_n685), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n599), .A2(G179), .A3(new_n532), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n480), .A2(new_n615), .A3(new_n496), .A4(new_n539), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n717), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n573), .B(G179), .C1(new_n582), .C2(new_n583), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n721), .A3(KEYINPUT30), .A4(new_n532), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n651), .B2(new_n611), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n605), .A2(new_n501), .A3(new_n540), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n725), .B2(new_n684), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n712), .B1(new_n714), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n684), .B1(new_n664), .B2(new_n674), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n711), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n705), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n274), .B1(new_n678), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n701), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n253), .A2(new_n468), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n241), .A2(G45), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n397), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n700), .B1(G355), .B2(new_n291), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n744), .A2(new_n745), .B1(G116), .B2(new_n700), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n238), .B1(G20), .B2(new_n311), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n741), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n749), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n239), .A2(G190), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n429), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n291), .B1(new_n758), .B2(G283), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n755), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G329), .ZN(new_n763));
  NAND3_X1  g0563(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT99), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT99), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(new_n304), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(KEYINPUT33), .B(G317), .Z(new_n768));
  OAI211_X1 g0568(.A(new_n759), .B(new_n763), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n765), .A2(G190), .A3(new_n766), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n239), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n770), .A2(new_n771), .B1(new_n773), .B2(new_n530), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT102), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n769), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n239), .A2(new_n304), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n756), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G303), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n351), .A2(G200), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n754), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n778), .B(new_n782), .C1(new_n783), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n779), .A2(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G322), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT103), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n781), .A2(G87), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n388), .A2(new_n389), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(new_n788), .B2(new_n793), .C1(new_n767), .C2(new_n202), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G107), .B2(new_n758), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n785), .A2(KEYINPUT98), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n785), .A2(KEYINPUT98), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n770), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n798), .A2(G77), .B1(G50), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n773), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G97), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n761), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n803), .A2(new_n291), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n791), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n750), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n752), .B1(new_n693), .B2(new_n753), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n693), .A2(G330), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n694), .B2(KEYINPUT97), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n693), .A2(KEYINPUT97), .A3(G330), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n813), .A2(new_n741), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n365), .A2(new_n684), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n432), .B2(new_n433), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n366), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n366), .A2(new_n684), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n732), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(new_n731), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n741), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n758), .A2(G68), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n397), .B1(new_n781), .B2(G50), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(new_n793), .C2(new_n773), .ZN(new_n831));
  INV_X1    g0631(.A(new_n767), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G150), .B1(G143), .B2(new_n789), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(new_n798), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n770), .C1(new_n835), .C2(new_n804), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT105), .B(KEYINPUT34), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n831), .B(new_n838), .C1(G132), .C2(new_n762), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n291), .B1(new_n798), .B2(G116), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n758), .A2(G87), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n802), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n762), .A2(G311), .B1(new_n799), .B2(G303), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n767), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n788), .A2(new_n530), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n780), .A2(new_n225), .ZN(new_n847));
  NOR4_X1   g0647(.A1(new_n842), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n750), .B1(new_n839), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n825), .A2(new_n747), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n750), .A2(new_n747), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n231), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n850), .A3(new_n740), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n828), .A2(new_n853), .ZN(G384));
  INV_X1    g0654(.A(KEYINPUT110), .ZN(new_n855));
  INV_X1    g0655(.A(new_n728), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n726), .C1(new_n644), .C2(new_n684), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n344), .A2(KEYINPUT107), .A3(new_n684), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n344), .A2(new_n684), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT107), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n345), .A2(new_n430), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n332), .A2(new_n344), .A3(new_n684), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n825), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n387), .A2(new_n407), .A3(new_n413), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n407), .A2(new_n413), .B1(new_n421), .B2(new_n682), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n405), .A2(new_n406), .A3(new_n273), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n413), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n422), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n682), .B1(new_n869), .B2(new_n413), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n874), .A3(new_n414), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n868), .B1(KEYINPUT37), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n426), .A2(KEYINPUT108), .A3(new_n873), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT108), .B1(new_n426), .B2(new_n873), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n877), .B(KEYINPUT38), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n865), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n855), .B1(new_n884), .B2(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n862), .A2(new_n863), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n366), .A2(new_n684), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n366), .B2(new_n822), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n714), .B2(new_n729), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n423), .A2(new_n425), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n873), .B1(new_n891), .B2(new_n647), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n426), .A2(KEYINPUT108), .A3(new_n873), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n896), .B2(new_n877), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n882), .B(new_n876), .C1(new_n894), .C2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n890), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(KEYINPUT110), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n867), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n414), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n866), .B2(new_n867), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT109), .ZN(new_n908));
  INV_X1    g0708(.A(new_n682), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n426), .A2(new_n418), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT109), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n882), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(new_n880), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n857), .A2(KEYINPUT40), .A3(new_n864), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT111), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n880), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT111), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n918), .A2(new_n890), .A3(new_n919), .A4(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n902), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n435), .A2(new_n857), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G330), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n883), .A2(KEYINPUT39), .A3(new_n880), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n345), .A2(new_n684), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n891), .A2(new_n682), .ZN(new_n932));
  INV_X1    g0732(.A(new_n674), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n685), .B(new_n888), .C1(new_n933), .C2(new_n663), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n883), .A2(new_n880), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n938), .A3(new_n886), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n436), .B1(new_n734), .B2(new_n711), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n650), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n925), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n274), .B2(new_n678), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n585), .B1(new_n442), .B2(KEYINPUT35), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(new_n240), .C1(KEYINPUT35), .C2(new_n442), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n241), .A2(G77), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n392), .A2(new_n394), .ZN(new_n950));
  INV_X1    g0750(.A(new_n207), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n949), .A2(new_n950), .B1(new_n202), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(G1), .A3(new_n214), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n945), .A2(new_n948), .A3(new_n953), .ZN(G367));
  NOR2_X1   g0754(.A1(new_n696), .A2(new_n520), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT42), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n642), .B(new_n500), .C1(new_n641), .C2(new_n685), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n666), .A2(new_n685), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(new_n560), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n685), .B1(new_n960), .B2(new_n671), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n630), .A2(new_n632), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n684), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n659), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n654), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n956), .A2(new_n961), .B1(KEYINPUT43), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n959), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n695), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n701), .B(KEYINPUT41), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n690), .A2(new_n694), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n975), .A2(new_n695), .A3(new_n696), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n977), .A2(new_n735), .A3(KEYINPUT113), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n976), .A2(new_n731), .A3(new_n711), .A4(new_n734), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT113), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n570), .A2(new_n687), .B1(new_n560), .B2(new_n685), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n959), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT112), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n984), .A3(new_n959), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n988), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT114), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n695), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n695), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT114), .ZN(new_n994));
  INV_X1    g0794(.A(new_n981), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n970), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n990), .A2(new_n992), .A3(new_n994), .A4(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI211_X1 g0800(.A(KEYINPUT114), .B(new_n993), .C1(new_n990), .C2(new_n998), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n978), .B(new_n980), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n974), .B1(new_n1002), .B2(new_n736), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n972), .B1(new_n1003), .B2(new_n739), .ZN(new_n1004));
  INV_X1    g0804(.A(G317), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n761), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT46), .B1(new_n781), .B2(G116), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G107), .B2(new_n801), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n397), .C1(new_n530), .C2(new_n767), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1006), .B(new_n1009), .C1(G283), .C2(new_n798), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n799), .A2(G311), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n758), .A2(G97), .B1(G303), .B2(new_n789), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n799), .A2(G143), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n758), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n835), .A2(new_n207), .B1(new_n231), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G159), .B2(new_n832), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n397), .B1(new_n789), .B2(G150), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n801), .A2(G68), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n761), .A2(new_n834), .B1(new_n793), .B2(new_n780), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT115), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1014), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n750), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n964), .A2(new_n749), .A3(new_n965), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n700), .A2(new_n291), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n751), .B1(new_n216), .B2(new_n359), .C1(new_n249), .C2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n740), .A3(new_n1027), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1004), .A2(new_n1031), .ZN(G387));
  AOI22_X1  g0832(.A1(new_n798), .A2(G303), .B1(G322), .B2(new_n799), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n783), .B2(new_n767), .C1(new_n1005), .C2(new_n788), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT48), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n844), .B2(new_n773), .C1(new_n530), .C2(new_n780), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n397), .B1(new_n771), .B2(new_n761), .C1(new_n1016), .C2(new_n585), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n780), .A2(new_n231), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n773), .A2(new_n359), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n832), .B2(new_n263), .ZN(new_n1043));
  INV_X1    g0843(.A(G150), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n761), .C1(new_n804), .C2(new_n770), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1041), .B(new_n1045), .C1(G50), .C2(new_n789), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n291), .C1(new_n202), .C2(new_n786), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G97), .B2(new_n758), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n750), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n246), .A2(new_n468), .A3(new_n291), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n356), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(G68), .A2(G77), .ZN(new_n1052));
  OAI21_X1  g0852(.A(KEYINPUT50), .B1(new_n356), .B2(G50), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n468), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n702), .B1(new_n1054), .B2(new_n397), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n216), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n751), .C1(new_n225), .C2(new_n216), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n686), .A2(new_n689), .A3(new_n749), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1049), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1059), .A2(new_n740), .B1(new_n739), .B2(new_n976), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n977), .A2(new_n735), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n701), .A3(new_n979), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(G393));
  NAND3_X1  g0863(.A1(new_n990), .A2(new_n994), .A3(new_n998), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n992), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n979), .A3(new_n999), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1002), .A2(new_n701), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT117), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT117), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1066), .A2(new_n1070), .A3(new_n999), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n739), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n959), .A2(new_n753), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT118), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n770), .A2(new_n1005), .B1(new_n783), .B2(new_n788), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  INV_X1    g0876(.A(G303), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n397), .C1(new_n1077), .C2(new_n767), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G283), .B2(new_n781), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n801), .A2(G116), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n762), .A2(G322), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n758), .A2(G107), .B1(G294), .B2(new_n785), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n801), .A2(G77), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n202), .B2(new_n780), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n397), .B(new_n1085), .C1(new_n798), .C2(new_n357), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n762), .A2(G143), .B1(new_n832), .B2(new_n951), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n770), .A2(new_n1044), .B1(new_n804), .B2(new_n788), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1086), .A2(new_n841), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n810), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n751), .B1(new_n221), .B2(new_n216), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n256), .B2(new_n1028), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1091), .A2(new_n741), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1073), .A2(KEYINPUT118), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1074), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1068), .A2(new_n1072), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  AND4_X1   g0898(.A1(G330), .A2(new_n857), .A3(new_n888), .A4(new_n886), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n937), .A2(new_n886), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n930), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(new_n927), .B2(new_n928), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n918), .A2(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n709), .A2(new_n685), .A3(new_n823), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n824), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1105), .B2(new_n886), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1099), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1106), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1099), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n930), .B1(new_n937), .B2(new_n886), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n1109), .C1(new_n929), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1112), .A2(new_n738), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n851), .A2(new_n262), .A3(new_n261), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n929), .A2(new_n748), .ZN(new_n1115));
  INV_X1    g0915(.A(G132), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n788), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n780), .A2(new_n1044), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n291), .C1(new_n1120), .C2(new_n770), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G137), .B2(new_n832), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n804), .B2(new_n773), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI211_X1 g0924(.A(new_n1117), .B(new_n1123), .C1(new_n798), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n761), .C1(new_n207), .C2(new_n1016), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n798), .A2(G97), .B1(G283), .B2(new_n799), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n225), .B2(new_n767), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n762), .A2(G294), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1131), .A2(new_n829), .A3(new_n792), .A4(new_n1084), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n291), .B(new_n1132), .C1(G116), .C2(new_n789), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n810), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1115), .A2(new_n741), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1113), .B1(new_n1114), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n886), .B1(new_n730), .B2(new_n888), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n937), .B1(new_n1138), .B2(new_n1099), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n1138), .A2(new_n1105), .A3(new_n1099), .ZN(new_n1142));
  OAI211_X1 g0942(.A(KEYINPUT119), .B(new_n937), .C1(new_n1138), .C2(new_n1099), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n923), .A2(new_n712), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n941), .A2(new_n1145), .A3(new_n650), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1112), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1107), .A2(new_n1111), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n701), .A3(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(KEYINPUT120), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(KEYINPUT120), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1137), .B1(new_n1151), .B2(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(KEYINPUT123), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n855), .B(KEYINPUT40), .C1(new_n938), .C2(new_n890), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT110), .B1(new_n899), .B2(new_n900), .ZN(new_n1156));
  OAI211_X1 g0956(.A(G330), .B(new_n921), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n309), .B2(new_n313), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n309), .A2(new_n313), .A3(new_n1159), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1161), .A2(new_n284), .A3(new_n909), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n284), .A2(new_n909), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1162), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n1160), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1157), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n940), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1167), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n902), .A2(G330), .A3(new_n921), .A4(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1169), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1154), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT123), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1149), .A2(new_n1146), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n940), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1175), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(KEYINPUT57), .A3(new_n1178), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n701), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1167), .A2(new_n747), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n229), .B1(new_n372), .B2(G41), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n770), .A2(new_n1126), .B1(new_n786), .B2(new_n834), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n781), .A2(new_n1124), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT122), .Z(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(G150), .C2(new_n801), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n1120), .B2(new_n788), .C1(new_n1116), .C2(new_n767), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n758), .A2(G159), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n762), .B2(G124), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1193), .A2(new_n529), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1187), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1041), .B1(G107), .B2(new_n789), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n844), .B2(new_n761), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n291), .A2(G41), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1020), .B(new_n1201), .C1(new_n585), .C2(new_n770), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n786), .A2(new_n359), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1200), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n758), .B1(new_n389), .B2(new_n388), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n221), .C2(new_n767), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT58), .Z(new_n1207));
  OAI21_X1  g1007(.A(new_n750), .B1(new_n1198), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n851), .A2(new_n207), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1186), .A2(new_n740), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1177), .B2(new_n739), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1185), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(G375));
  INV_X1    g1015(.A(new_n1144), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1146), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n973), .A3(new_n1147), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n761), .A2(new_n1077), .B1(new_n770), .B2(new_n530), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1042), .B(new_n1220), .C1(G116), .C2(new_n832), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n397), .B1(new_n788), .B2(new_n844), .C1(new_n221), .C2(new_n780), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G77), .B2(new_n758), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(new_n225), .C2(new_n835), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n801), .A2(G50), .B1(new_n781), .B2(G159), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1044), .B2(new_n786), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1205), .A2(new_n291), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(G128), .C2(new_n762), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT124), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n832), .A2(new_n1124), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n834), .C2(new_n788), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n770), .A2(new_n1116), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n750), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n740), .C1(new_n748), .C2(new_n886), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n202), .B2(new_n851), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1144), .B2(new_n739), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1219), .A2(new_n1237), .ZN(G381));
  AND2_X1   g1038(.A1(new_n1137), .A2(new_n1150), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1214), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  INV_X1    g1041(.A(G381), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1097), .A2(new_n1004), .A3(new_n1031), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1060), .A2(new_n819), .A3(new_n1062), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n683), .A2(G213), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT125), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1240), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G378), .B(new_n1212), .C1(new_n1179), .C2(new_n1184), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT123), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1176), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n973), .B(new_n1178), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1211), .B1(new_n1182), .B2(new_n739), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1239), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1252), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1218), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1216), .A2(new_n1217), .A3(KEYINPUT60), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n701), .A4(new_n1147), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(G384), .A3(new_n1237), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G384), .B1(new_n1263), .B2(new_n1237), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G2897), .B(new_n1248), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1266), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1251), .A2(G2897), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1264), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT63), .B1(new_n1259), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1259), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1097), .A2(new_n1004), .A3(new_n1031), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1072), .A2(new_n1096), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1004), .A2(new_n1031), .B1(new_n1277), .B2(new_n1068), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1244), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT126), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1282), .A3(new_n1244), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1276), .A2(new_n1278), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1284), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1243), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1248), .B1(new_n1252), .B2(new_n1258), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1273), .A2(KEYINPUT63), .ZN(new_n1291));
  AOI211_X1 g1091(.A(KEYINPUT61), .B(new_n1289), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1275), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1259), .A2(new_n1294), .A3(new_n1273), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1273), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1296), .B2(KEYINPUT62), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT62), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1290), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1289), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(G405));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1289), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1289), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT127), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1239), .B1(new_n1185), .B2(new_n1213), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1296), .A3(new_n1252), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1296), .B1(new_n1306), .B2(new_n1252), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1303), .B(new_n1305), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1309), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(KEYINPUT127), .A3(new_n1304), .A4(new_n1307), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(G402));
endmodule


