//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n199), .A2(KEYINPUT64), .A3(G146), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT64), .B1(new_n199), .B2(G146), .ZN(new_n201));
  OAI211_X1 g015(.A(G128), .B(new_n198), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n199), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n197), .B2(G143), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT64), .A3(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n202), .A2(KEYINPUT1), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT80), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT79), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n216), .B(new_n218), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n212), .A2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n213), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n214), .A2(new_n215), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n218), .B2(new_n224), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n210), .A2(new_n226), .A3(KEYINPUT82), .A4(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n214), .A2(new_n225), .A3(new_n223), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G101), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(KEYINPUT81), .A3(new_n236), .A4(G101), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n199), .A2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n198), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n245), .B(new_n198), .C1(new_n200), .C2(new_n201), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n207), .A2(new_n250), .A3(new_n245), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n235), .A2(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n241), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n226), .A2(new_n227), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n209), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n243), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n244), .B2(new_n209), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n207), .A2(new_n262), .A3(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n234), .A2(new_n255), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G137), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT67), .A2(G137), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT67), .A2(G137), .ZN(new_n270));
  OAI211_X1 g084(.A(KEYINPUT11), .B(G134), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT66), .B(new_n272), .C1(new_n267), .C2(G137), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G134), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT66), .B1(new_n276), .B2(new_n272), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n268), .B(new_n271), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G131), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n272), .B1(new_n267), .B2(G137), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n273), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n268), .A4(new_n271), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT85), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n266), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n234), .A2(new_n255), .A3(new_n287), .A4(new_n265), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n196), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n286), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n234), .A2(new_n255), .A3(new_n292), .A4(new_n265), .ZN(new_n293));
  INV_X1    g107(.A(new_n264), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n230), .A2(new_n231), .B1(new_n294), .B2(new_n256), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT12), .B1(new_n295), .B2(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n256), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n232), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n286), .ZN(new_n300));
  AND4_X1   g114(.A1(new_n196), .A2(new_n293), .A3(new_n296), .A4(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n191), .B(new_n192), .C1(new_n291), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT86), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n289), .A2(new_n290), .ZN(new_n304));
  INV_X1    g118(.A(new_n196), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n293), .A2(new_n300), .A3(new_n196), .A4(new_n296), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n191), .A4(new_n192), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n296), .A3(new_n300), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n196), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n293), .A2(new_n300), .A3(KEYINPUT84), .A4(new_n296), .ZN(new_n315));
  INV_X1    g129(.A(new_n304), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n196), .ZN(new_n317));
  OAI21_X1  g131(.A(G469), .B1(new_n317), .B2(G902), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n190), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n286), .A2(new_n252), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n269), .A2(new_n270), .A3(G134), .ZN(new_n322));
  INV_X1    g136(.A(new_n276), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n264), .A2(new_n285), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT73), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  INV_X1    g142(.A(G116), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G116), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n329), .A2(G119), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT70), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT2), .B(G113), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT70), .ZN(new_n337));
  INV_X1    g151(.A(new_n334), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT69), .B(G116), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n328), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n338), .B1(new_n339), .B2(new_n328), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n342), .A2(new_n336), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n341), .B2(new_n343), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n321), .A2(new_n349), .A3(new_n325), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n327), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n326), .A2(new_n347), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n321), .B(new_n325), .C1(new_n345), .C2(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n355));
  AOI22_X1  g169(.A1(new_n320), .A2(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(G101), .ZN(new_n358));
  NOR2_X1   g172(.A1(G237), .A2(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G210), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT74), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n321), .A2(new_n363), .A3(new_n325), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n321), .B2(new_n325), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n347), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n353), .A3(new_n361), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT31), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n366), .A2(KEYINPUT31), .A3(new_n353), .A4(new_n361), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n351), .A2(new_n320), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n354), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n375));
  INV_X1    g189(.A(new_n361), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n362), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G472), .A2(G902), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n361), .B1(new_n366), .B2(new_n353), .ZN(new_n384));
  AOI211_X1 g198(.A(KEYINPUT29), .B(new_n384), .C1(new_n361), .C2(new_n356), .ZN(new_n385));
  INV_X1    g199(.A(new_n354), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n372), .B1(new_n320), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n361), .A2(KEYINPUT29), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n192), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G472), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(G234), .A2(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G952), .A3(new_n194), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT21), .B(G898), .Z(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(G902), .A3(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n217), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n194), .A3(G214), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n199), .ZN(new_n410));
  AOI21_X1  g224(.A(G143), .B1(new_n359), .B2(G214), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n199), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n359), .A2(G143), .A3(G214), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n413), .A2(KEYINPUT18), .A3(G131), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G125), .B(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n197), .ZN(new_n418));
  INV_X1    g232(.A(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G125), .ZN(new_n420));
  INV_X1    g234(.A(G125), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G140), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT77), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n421), .A2(KEYINPUT77), .A3(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n418), .B1(new_n425), .B2(new_n197), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT16), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n423), .B2(new_n424), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n420), .A2(KEYINPUT16), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n197), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n421), .A2(KEYINPUT77), .A3(G140), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n417), .B2(KEYINPUT77), .ZN(new_n435));
  OAI211_X1 g249(.A(G146), .B(new_n433), .C1(new_n435), .C2(new_n429), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT78), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n430), .A2(new_n431), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(G146), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G131), .B1(new_n410), .B2(new_n411), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n413), .A2(new_n284), .A3(new_n414), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT17), .ZN(new_n445));
  MUX2_X1   g259(.A(new_n442), .B(new_n444), .S(new_n445), .Z(new_n446));
  AOI211_X1 g260(.A(new_n406), .B(new_n428), .C1(new_n441), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n417), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n425), .B2(new_n449), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n436), .B(new_n444), .C1(new_n451), .C2(G146), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n427), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n453), .B2(new_n406), .ZN(new_n454));
  AOI211_X1 g268(.A(KEYINPUT91), .B(new_n405), .C1(new_n452), .C2(new_n427), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n447), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G475), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n192), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n454), .ZN(new_n460));
  INV_X1    g274(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n441), .A2(new_n446), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n405), .A3(new_n427), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n464), .A2(new_n465), .A3(new_n457), .A4(new_n192), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n405), .B1(new_n462), .B2(new_n427), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n192), .B1(new_n468), .B2(new_n447), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT92), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(new_n192), .C1(new_n468), .C2(new_n447), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(G475), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n474));
  INV_X1    g288(.A(G122), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n330), .B2(new_n332), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n329), .A2(G122), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT93), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n479));
  INV_X1    g293(.A(new_n477), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(new_n480), .C1(new_n339), .C2(new_n475), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n478), .A2(new_n212), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n212), .B1(new_n478), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n481), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G107), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n478), .A2(new_n212), .A3(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(KEYINPUT94), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n199), .A2(G128), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n208), .A2(G143), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(new_n267), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT13), .B1(new_n199), .B2(G128), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT95), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT13), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n494), .B(new_n490), .C1(new_n495), .C2(new_n489), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n492), .B1(new_n496), .B2(G134), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n484), .A2(new_n488), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n476), .A2(KEYINPUT14), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n330), .A2(new_n332), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G122), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n480), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n499), .B(G107), .C1(new_n502), .C2(KEYINPUT14), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n491), .A2(new_n267), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n503), .B(new_n487), .C1(new_n492), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G217), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n188), .A2(new_n507), .A3(G953), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n498), .A2(new_n505), .A3(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n192), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n512), .B(new_n192), .C1(KEYINPUT15), .C2(new_n514), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n467), .A2(new_n473), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n346), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n241), .A2(new_n519), .A3(new_n520), .A4(new_n254), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n335), .B2(new_n340), .ZN(new_n523));
  OAI21_X1  g337(.A(G113), .B1(new_n338), .B2(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n343), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n525), .A2(new_n256), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT6), .ZN(new_n529));
  XOR2_X1   g343(.A(G110), .B(G122), .Z(new_n530));
  NAND4_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n294), .A2(new_n421), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n421), .B2(new_n252), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n194), .A2(G224), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT88), .Z(new_n535));
  XOR2_X1   g349(.A(new_n533), .B(new_n535), .Z(new_n536));
  INV_X1    g350(.A(new_n530), .ZN(new_n537));
  AOI211_X1 g351(.A(KEYINPUT87), .B(new_n537), .C1(new_n521), .C2(new_n526), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n521), .A2(new_n537), .A3(new_n526), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT6), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n531), .B(new_n536), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n533), .B(new_n542), .Z(new_n543));
  OR2_X1    g357(.A1(new_n525), .A2(new_n257), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n530), .B(KEYINPUT8), .Z(new_n545));
  NOR2_X1   g359(.A1(new_n342), .A2(new_n522), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n343), .B1(new_n546), .B2(new_n524), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n257), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT89), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n544), .A2(new_n551), .A3(new_n545), .A4(new_n548), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n543), .A2(new_n539), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n541), .A2(new_n192), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G210), .B1(G237), .B2(G902), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT90), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n541), .A2(new_n553), .A3(new_n192), .A4(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n403), .B(new_n518), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n328), .A2(G128), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(G119), .B2(new_n208), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  INV_X1    g379(.A(KEYINPUT23), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(G119), .B2(new_n208), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n328), .A2(KEYINPUT23), .A3(G128), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n564), .A2(new_n565), .B1(G110), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n436), .A3(new_n418), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(new_n565), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n437), .A2(new_n572), .A3(new_n440), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(G110), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT76), .Z(new_n575));
  OAI21_X1  g389(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT22), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G137), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n576), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n192), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT25), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n507), .B1(G234), .B2(new_n192), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n584), .A3(new_n192), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n583), .A2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n319), .A2(new_n391), .A3(new_n560), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  INV_X1    g405(.A(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n378), .B2(new_n192), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n379), .B2(new_n378), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n319), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n511), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n512), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n510), .B(new_n511), .C1(new_n598), .C2(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n514), .A2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT97), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n513), .A2(new_n514), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n602), .A2(new_n607), .A3(new_n603), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n467), .A2(new_n473), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n554), .A2(new_n555), .ZN(new_n612));
  INV_X1    g426(.A(new_n555), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n541), .A2(new_n553), .A3(new_n192), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n402), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n596), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND2_X1  g433(.A1(new_n516), .A2(new_n517), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n466), .A2(KEYINPUT98), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n459), .A2(KEYINPUT98), .A3(new_n466), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n473), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n596), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  INV_X1    g441(.A(new_n579), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n576), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n587), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n586), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n319), .A2(new_n594), .A3(new_n560), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT99), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT37), .B(G110), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  NAND3_X1  g450(.A1(new_n612), .A2(new_n400), .A3(new_n614), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n319), .A2(new_n391), .A3(new_n632), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n393), .B(KEYINPUT100), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n398), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n623), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n208), .ZN(G30));
  AND2_X1   g460(.A1(new_n557), .A2(new_n559), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT38), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n366), .A2(new_n353), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n361), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n192), .C1(new_n361), .C2(new_n354), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G472), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n382), .A2(new_n652), .A3(new_n383), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n467), .A2(new_n473), .B1(new_n516), .B2(new_n517), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n400), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n632), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n642), .B(KEYINPUT39), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n319), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT40), .B1(new_n319), .B2(new_n660), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n199), .ZN(G45));
  INV_X1    g481(.A(new_n642), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n609), .A2(new_n610), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n639), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n197), .ZN(G48));
  AND2_X1   g485(.A1(new_n391), .A2(new_n589), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n306), .B2(new_n307), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n191), .B1(new_n674), .B2(KEYINPUT101), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n192), .B1(new_n291), .B2(new_n301), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n675), .A2(new_n678), .B1(new_n303), .B2(new_n310), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n673), .B1(new_n679), .B2(new_n189), .ZN(new_n680));
  OAI211_X1 g494(.A(KEYINPUT101), .B(new_n192), .C1(new_n291), .C2(new_n301), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n678), .A2(G469), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n311), .A2(new_n682), .A3(new_n189), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n672), .B(new_n616), .C1(new_n680), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  OAI211_X1 g501(.A(new_n672), .B(new_n624), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n683), .B2(new_n637), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n679), .A2(new_n691), .A3(new_n638), .A4(new_n189), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n518), .ZN(new_n694));
  INV_X1    g508(.A(new_n399), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n391), .A2(new_n694), .A3(new_n695), .A4(new_n632), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NAND2_X1  g512(.A1(new_n387), .A2(new_n376), .ZN(new_n699));
  AOI211_X1 g513(.A(G472), .B(G902), .C1(new_n699), .C2(new_n371), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n593), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n589), .A3(new_n695), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n400), .A2(new_n612), .A3(new_n614), .A4(new_n656), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n702), .B(new_n703), .C1(new_n680), .C2(new_n684), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  INV_X1    g519(.A(new_n669), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n658), .A2(new_n593), .A3(new_n700), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n692), .B2(new_n690), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n421), .ZN(G27));
  NAND2_X1  g524(.A1(G469), .A2(G902), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT104), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n289), .A2(new_n290), .A3(new_n196), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n289), .A2(new_n715), .A3(new_n290), .A4(new_n196), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n314), .A2(new_n315), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(G469), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n309), .B1(new_n674), .B2(new_n191), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n302), .A2(KEYINPUT86), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n712), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n722), .A2(KEYINPUT42), .A3(new_n189), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n557), .A2(new_n559), .A3(new_n400), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n669), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n378), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n383), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n382), .A3(new_n390), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n723), .A2(new_n589), .A3(new_n726), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n391), .A2(new_n589), .A3(new_n724), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n722), .A2(new_n189), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n733), .A2(new_n669), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n732), .B1(new_n735), .B2(KEYINPUT42), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  INV_X1    g551(.A(new_n733), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n714), .A2(new_n716), .B1(new_n314), .B2(new_n315), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n303), .A2(new_n310), .B1(new_n739), .B2(G469), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n190), .B1(new_n740), .B2(new_n712), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n644), .A2(KEYINPUT107), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n644), .A2(KEYINPUT107), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n741), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n610), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT43), .A3(new_n609), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(KEYINPUT111), .A3(KEYINPUT43), .A4(new_n609), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n752));
  INV_X1    g566(.A(new_n609), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(new_n610), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n594), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(KEYINPUT44), .A3(new_n756), .A4(new_n632), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n632), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n725), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n739), .A2(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n718), .A2(new_n713), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n764), .A3(G469), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n712), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(new_n767), .B1(new_n310), .B2(new_n303), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n190), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT108), .A3(new_n660), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT108), .B1(new_n770), .B2(new_n660), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n757), .B(new_n760), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  INV_X1    g589(.A(new_n726), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n768), .A2(new_n769), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n777), .B1(new_n778), .B2(new_n190), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n391), .A2(new_n589), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(new_n190), .A2(new_n401), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n747), .A2(new_n589), .A3(new_n609), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT112), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n679), .B(KEYINPUT49), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n648), .A3(new_n654), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n725), .A2(new_n683), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n755), .A2(new_n790), .A3(new_n640), .A4(new_n707), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n683), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n648), .A2(new_n401), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n701), .A2(new_n589), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n640), .A3(new_n796), .A4(new_n755), .ZN(new_n797));
  OR2_X1    g611(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n589), .A2(new_n790), .A3(new_n394), .A4(new_n654), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n467), .A3(new_n473), .A4(new_n753), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n793), .A2(new_n799), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n679), .A2(new_n190), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n779), .A2(new_n780), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n755), .A2(new_n640), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(new_n796), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n724), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT51), .B1(new_n804), .B2(KEYINPUT119), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n815));
  INV_X1    g629(.A(new_n811), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n804), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n802), .A2(new_n610), .A3(new_n609), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n809), .A2(new_n589), .A3(new_n731), .A4(new_n790), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT48), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n194), .A2(G952), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n810), .B2(new_n693), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n706), .A2(new_n707), .A3(new_n722), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n621), .A2(new_n622), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n311), .B2(new_n318), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n473), .A2(new_n516), .A3(new_n517), .A4(new_n668), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n391), .A3(new_n632), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n647), .A3(new_n785), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n736), .A2(new_n832), .A3(new_n744), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n697), .A2(new_n685), .A3(new_n688), .A4(new_n704), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n647), .A2(new_n403), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n605), .A2(new_n610), .A3(new_n606), .A4(new_n608), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(KEYINPUT113), .A3(new_n518), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT113), .B1(new_n609), .B2(new_n610), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n590), .B(new_n633), .C1(new_n839), .C2(new_n595), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n632), .A2(new_n642), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT32), .B1(new_n378), .B2(new_n379), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n727), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n652), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n703), .A4(new_n741), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n653), .A2(new_n843), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n722), .A2(new_n703), .A3(new_n189), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT114), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n693), .A2(new_n706), .A3(new_n707), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n319), .A2(new_n638), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n658), .B1(new_n846), .B2(new_n390), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(new_n856), .C1(new_n643), .C2(new_n706), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT52), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n639), .B1(new_n644), .B2(new_n669), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n709), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n853), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n825), .B1(new_n842), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n862), .B1(new_n861), .B2(new_n853), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n862), .A2(new_n853), .A3(new_n854), .A4(new_n857), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n391), .A2(new_n589), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n679), .A2(new_n673), .A3(new_n189), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n872), .A2(new_n616), .B1(new_n693), .B2(new_n696), .ZN(new_n873));
  INV_X1    g687(.A(new_n840), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n688), .A4(new_n704), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n736), .A2(new_n832), .A3(new_n744), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n865), .A2(new_n878), .A3(KEYINPUT54), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT54), .B1(new_n865), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n824), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n842), .A2(new_n864), .A3(new_n825), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n868), .B2(new_n877), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n865), .A2(new_n878), .A3(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(KEYINPUT115), .A3(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n814), .B(new_n823), .C1(new_n881), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n789), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n194), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n192), .B1(new_n865), .B2(new_n878), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n893), .B2(G210), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n894), .B2(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n531), .B1(new_n538), .B2(new_n540), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n536), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(KEYINPUT120), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n895), .B1(new_n900), .B2(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n712), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n712), .A2(new_n904), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n885), .A2(new_n886), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n308), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n893), .A2(G469), .A3(new_n764), .A4(new_n761), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n891), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n911), .A2(G475), .A3(new_n464), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n464), .B1(new_n911), .B2(G475), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n891), .ZN(G60));
  INV_X1    g728(.A(new_n602), .ZN(new_n915));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  NOR4_X1   g731(.A1(new_n879), .A2(new_n880), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n881), .A2(new_n887), .A3(new_n919), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n891), .B(new_n918), .C1(new_n920), .C2(new_n915), .ZN(G63));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n865), .B2(new_n878), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n630), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n892), .B1(new_n925), .B2(new_n580), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n922), .B(KEYINPUT61), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n926), .B(new_n892), .C1(new_n580), .C2(new_n925), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT61), .B1(new_n931), .B2(new_n922), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(G66));
  INV_X1    g747(.A(G224), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n396), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n875), .B(KEYINPUT123), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n897), .B1(G898), .B2(new_n194), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NOR2_X1   g753(.A1(new_n364), .A2(new_n365), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(new_n451), .Z(new_n941));
  AND2_X1   g755(.A1(new_n760), .A2(new_n757), .ZN(new_n942));
  INV_X1    g756(.A(new_n773), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n771), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n942), .A2(new_n944), .B1(new_n781), .B2(new_n782), .ZN(new_n945));
  INV_X1    g759(.A(new_n838), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n836), .A2(KEYINPUT113), .A3(new_n518), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n319), .B(new_n660), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n733), .B(new_n950), .C1(new_n949), .C2(new_n948), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  INV_X1    g766(.A(new_n861), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n666), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n861), .B(KEYINPUT62), .C1(new_n665), .C2(new_n657), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n945), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n941), .B1(new_n957), .B2(G953), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n194), .A2(G900), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n736), .A2(new_n744), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n731), .A2(new_n589), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n943), .B2(new_n771), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(new_n703), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n774), .A2(KEYINPUT126), .A3(new_n861), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT126), .B1(new_n774), .B2(new_n861), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n783), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n194), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n958), .B1(new_n968), .B2(new_n941), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n958), .C1(new_n968), .C2(new_n941), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(G72));
  NAND3_X1  g788(.A1(new_n945), .A2(new_n936), .A3(new_n956), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  AOI21_X1  g791(.A(new_n650), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  INV_X1    g793(.A(new_n936), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n977), .B1(new_n967), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n649), .A2(new_n361), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n891), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n865), .A2(new_n878), .ZN(new_n984));
  INV_X1    g798(.A(new_n982), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n650), .A3(new_n977), .A4(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n979), .A2(new_n983), .A3(new_n986), .ZN(G57));
endmodule


