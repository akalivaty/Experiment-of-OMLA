//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G77), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G87), .A2(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT67), .Z(new_n225));
  AOI22_X1  g0025(.A1(new_n219), .A2(new_n225), .B1(G1), .B2(G20), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n211), .B(new_n227), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT69), .Z(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n260), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n266), .A2(G223), .B1(new_n215), .B2(new_n265), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n254), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n252), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n214), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n228), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n229), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT70), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n203), .A2(new_n229), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n280), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n213), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n280), .B1(new_n251), .B2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n278), .B(new_n295), .C1(G179), .C2(new_n276), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT71), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n214), .A2(new_n260), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n235), .A2(G1698), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n299), .B(new_n300), .C1(new_n263), .C2(new_n264), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n254), .B1(new_n303), .B2(new_n271), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n270), .A2(G238), .A3(new_n252), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n270), .B1(new_n301), .B2(new_n302), .ZN(new_n308));
  NOR4_X1   g0108(.A1(new_n308), .A2(KEYINPUT13), .A3(new_n305), .A4(new_n254), .ZN(new_n309));
  OAI21_X1  g0109(.A(G169), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT14), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n307), .A2(new_n309), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G179), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(G169), .C1(new_n307), .C2(new_n309), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G68), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G20), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n318), .B1(new_n282), .B2(new_n204), .C1(new_n285), .C2(new_n213), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n280), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT11), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(new_n321), .B1(G68), .B2(new_n293), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT76), .B1(new_n290), .B2(G68), .ZN(new_n324));
  XOR2_X1   g0124(.A(new_n324), .B(KEYINPUT12), .Z(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n304), .A2(new_n306), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(new_n309), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n326), .B1(new_n331), .B2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n312), .A2(G190), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n276), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n272), .B2(new_n275), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT75), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT10), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n295), .B(KEYINPUT9), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n340), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n297), .B(new_n335), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n347));
  INV_X1    g0147(.A(new_n281), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n291), .ZN(new_n349));
  INV_X1    g0149(.A(new_n293), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n257), .A2(new_n229), .A3(new_n258), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n258), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n317), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G58), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n317), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n358), .B2(new_n201), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n284), .A2(G159), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT16), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n265), .B2(new_n229), .ZN(new_n363));
  INV_X1    g0163(.A(new_n355), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  INV_X1    g0166(.A(new_n361), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n351), .B1(new_n369), .B2(new_n280), .ZN(new_n370));
  OR2_X1    g0170(.A1(G223), .A2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n214), .A2(G1698), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n372), .C1(new_n263), .C2(new_n264), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n271), .ZN(new_n376));
  INV_X1    g0176(.A(new_n273), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G232), .ZN(new_n378));
  INV_X1    g0178(.A(new_n254), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n376), .A2(G190), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n270), .B1(new_n373), .B2(new_n374), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n273), .A2(new_n235), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(new_n254), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n383), .B2(new_n338), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n347), .B1(new_n370), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n280), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n362), .B2(new_n368), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NOR4_X1   g0190(.A1(new_n388), .A2(new_n384), .A3(new_n351), .A4(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n376), .A2(G179), .A3(new_n378), .A4(new_n379), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n383), .B2(new_n277), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n393), .B1(new_n370), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(KEYINPUT18), .C1(new_n388), .C2(new_n351), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n215), .A2(G20), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n401), .B1(new_n285), .B2(new_n281), .C1(new_n402), .C2(new_n282), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT73), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(new_n280), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n403), .B2(new_n280), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n293), .A2(G77), .B1(new_n216), .B2(new_n291), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n266), .A2(G238), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n265), .A2(G107), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n259), .A2(new_n414), .A3(G232), .A4(new_n260), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n271), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n273), .A2(new_n217), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n417), .A2(G190), .A3(new_n379), .A4(new_n419), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n254), .B(new_n418), .C1(new_n416), .C2(new_n271), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n409), .B(new_n420), .C1(new_n338), .C2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n417), .A2(new_n423), .A3(new_n379), .A4(new_n419), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n403), .A2(new_n280), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT73), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n403), .A2(new_n404), .A3(new_n280), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n407), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n424), .B(new_n428), .C1(new_n421), .C2(G169), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n430), .B(KEYINPUT74), .Z(new_n431));
  NOR3_X1   g0231(.A1(new_n346), .A2(new_n400), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(KEYINPUT6), .A3(G97), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n222), .A2(new_n433), .ZN(new_n435));
  NOR2_X1   g0235(.A1(G97), .A2(G107), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n434), .B1(new_n437), .B2(KEYINPUT6), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n439));
  OAI21_X1  g0239(.A(G107), .B1(new_n363), .B2(new_n364), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n280), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n256), .A2(G1), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n228), .B(new_n279), .C1(new_n443), .C2(KEYINPUT78), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n251), .A2(KEYINPUT78), .A3(G33), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n290), .A2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n444), .A2(new_n446), .A3(KEYINPUT79), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT78), .B1(new_n251), .B2(G33), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n280), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n290), .A2(new_n445), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(G97), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n290), .A2(G97), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT80), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT79), .B1(new_n444), .B2(new_n446), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n451), .A3(new_n448), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n222), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT80), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n459), .A2(new_n460), .A3(new_n454), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n442), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n251), .A2(G45), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(G41), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT5), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n464), .A2(new_n466), .A3(new_n468), .A4(G274), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n251), .B(G45), .C1(new_n465), .C2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n467), .A2(KEYINPUT5), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n270), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(new_n223), .ZN(new_n473));
  OAI211_X1 g0273(.A(G244), .B(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT4), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n473), .B1(new_n480), .B2(new_n271), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G169), .ZN(new_n482));
  AOI211_X1 g0282(.A(G179), .B(new_n473), .C1(new_n480), .C2(new_n271), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n462), .A2(new_n484), .ZN(new_n485));
  OR2_X1    g0285(.A1(G238), .A2(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n217), .A2(G1698), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n487), .C1(new_n263), .C2(new_n264), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G116), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n270), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n270), .A2(G250), .A3(new_n463), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n464), .A2(G274), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n490), .A2(new_n493), .A3(G179), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT81), .ZN(new_n495));
  INV_X1    g0295(.A(new_n402), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n290), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n282), .B2(new_n222), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT82), .B(new_n498), .C1(new_n282), .C2(new_n222), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n229), .B1(new_n302), .B2(new_n498), .ZN(new_n503));
  INV_X1    g0303(.A(G87), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n436), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n229), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n501), .A2(new_n502), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n497), .B1(new_n508), .B2(new_n280), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n496), .B1(new_n447), .B2(new_n452), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n490), .A2(new_n493), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n509), .A2(new_n510), .B1(new_n512), .B2(new_n277), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n488), .A2(new_n489), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n271), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(G190), .A3(new_n492), .A4(new_n491), .ZN(new_n516));
  OAI21_X1  g0316(.A(G87), .B1(new_n447), .B2(new_n452), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n509), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(G200), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n495), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n453), .A2(KEYINPUT80), .A3(new_n455), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n460), .B1(new_n459), .B2(new_n454), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(new_n280), .B2(new_n441), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n481), .A2(new_n336), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G200), .B2(new_n481), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n485), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n528));
  OAI211_X1 g0328(.A(G257), .B(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n257), .A2(G303), .A3(new_n258), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n271), .ZN(new_n532));
  OAI211_X1 g0332(.A(G270), .B(new_n270), .C1(new_n470), .C2(new_n471), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n469), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n450), .A2(new_n451), .A3(G116), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n291), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n279), .A2(new_n228), .B1(G20), .B2(new_n536), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n478), .B(new_n229), .C1(G33), .C2(new_n222), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT20), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n535), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n534), .A2(G169), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n534), .A2(KEYINPUT21), .A3(new_n542), .A4(G169), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n532), .A2(new_n533), .A3(G179), .A4(new_n469), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n542), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n534), .A2(G200), .ZN(new_n551));
  INV_X1    g0351(.A(new_n542), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n336), .C2(new_n534), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n527), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n229), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT83), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(KEYINPUT22), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n556), .B(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n489), .A2(KEYINPUT84), .A3(G20), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT84), .B1(new_n489), .B2(G20), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT23), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n229), .B2(G107), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n433), .A2(KEYINPUT23), .A3(G20), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n561), .A2(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n559), .A2(new_n560), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n560), .B1(new_n559), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n280), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n447), .B2(new_n452), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n290), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n223), .A2(G1698), .ZN(new_n574));
  OAI221_X1 g0374(.A(new_n574), .B1(G250), .B2(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n270), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G264), .B(new_n270), .C1(new_n470), .C2(new_n471), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n469), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(G169), .ZN(new_n582));
  INV_X1    g0382(.A(new_n579), .ZN(new_n583));
  INV_X1    g0383(.A(new_n469), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT85), .B1(new_n585), .B2(new_n277), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n582), .B(new_n586), .C1(new_n423), .C2(new_n580), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n573), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(new_n336), .A3(new_n469), .A4(new_n579), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n585), .B2(G200), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n569), .A2(new_n590), .A3(new_n570), .A4(new_n572), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n594), .A3(new_n591), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n432), .A2(new_n555), .A3(new_n596), .ZN(G372));
  AND2_X1   g0397(.A1(new_n485), .A2(new_n526), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n491), .A2(new_n492), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n515), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n494), .B1(new_n509), .B2(new_n510), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n277), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n518), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n591), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n598), .A2(KEYINPUT88), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n485), .A2(new_n526), .A3(new_n591), .A4(new_n607), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n573), .B2(new_n587), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n609), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n481), .A2(new_n423), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G169), .B2(new_n481), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n523), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n520), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n605), .A2(new_n606), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n623), .A3(new_n607), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n432), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n361), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n280), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n351), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT18), .B1(new_n632), .B2(new_n395), .ZN(new_n633));
  INV_X1    g0433(.A(new_n398), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n370), .A2(new_n385), .A3(new_n389), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n388), .A2(new_n384), .A3(new_n351), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n347), .ZN(new_n638));
  INV_X1    g0438(.A(new_n429), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n334), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n640), .B2(new_n327), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n344), .A2(new_n345), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(new_n297), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n627), .A2(new_n643), .ZN(G369));
  XOR2_X1   g0444(.A(KEYINPUT89), .B(KEYINPUT27), .Z(new_n645));
  INV_X1    g0445(.A(G13), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n646), .A2(G1), .A3(G20), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n552), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n613), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n554), .B2(new_n654), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT90), .Z(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n588), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n573), .A2(new_n652), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n596), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n588), .A2(new_n652), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n550), .A2(new_n652), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n596), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n209), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n505), .A2(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n231), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n601), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n600), .B1(new_n491), .B2(new_n492), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n515), .B(KEYINPUT93), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n423), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT93), .B1(new_n602), .B2(new_n515), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n481), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n534), .A4(new_n580), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NOR4_X1   g0485(.A1(new_n577), .A2(new_n490), .A3(new_n583), .A4(new_n493), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n548), .B1(new_n686), .B2(KEYINPUT92), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n511), .A2(new_n578), .A3(new_n579), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n481), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n547), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT30), .A4(new_n481), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n684), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n652), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n698), .A3(new_n652), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n555), .A2(new_n593), .A3(new_n595), .A4(new_n653), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n676), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n619), .A2(new_n623), .A3(new_n520), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n622), .B(new_n703), .C1(new_n610), .C2(new_n614), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n623), .B1(new_n619), .B2(new_n607), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n653), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT94), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT94), .B(new_n653), .C1(new_n704), .C2(new_n705), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(new_n626), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n652), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n702), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n675), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR2_X1   g0516(.A1(new_n229), .A2(new_n336), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(new_n423), .A3(G200), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n229), .A2(G190), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n719), .A2(G322), .B1(G329), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n423), .A2(new_n338), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G326), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n265), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n338), .A2(G179), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n720), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n729), .B1(G283), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n229), .B1(new_n721), .B2(G190), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G294), .ZN(new_n736));
  INV_X1    g0536(.A(new_n720), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n737), .A2(new_n423), .A3(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n717), .A2(new_n730), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n738), .A2(G311), .B1(new_n740), .B2(G303), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n725), .A2(new_n720), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(KEYINPUT33), .A2(G317), .ZN(new_n744));
  AND2_X1   g0544(.A1(KEYINPUT33), .A2(G317), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n733), .A2(new_n736), .A3(new_n741), .A4(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n738), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT96), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n719), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n216), .B1(new_n357), .B2(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n753), .A2(KEYINPUT97), .B1(G68), .B2(new_n743), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n732), .A2(G107), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n734), .A2(new_n222), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G50), .A2(new_n727), .B1(new_n740), .B2(G87), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n754), .A2(new_n755), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G159), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n722), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT32), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n259), .B(new_n762), .C1(new_n753), .C2(KEYINPUT97), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n747), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT98), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n228), .B1(G20), .B2(new_n277), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n655), .B(new_n770), .C1(new_n554), .C2(new_n654), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n646), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G45), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n670), .A2(G1), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n668), .A2(new_n259), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n246), .B2(G45), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n231), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n259), .A2(new_n209), .ZN(new_n780));
  INV_X1    g0580(.A(G355), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n209), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT95), .Z(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n770), .A2(new_n766), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n767), .A2(new_n771), .A3(new_n775), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n658), .A2(new_n774), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n657), .A2(G330), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(G396));
  INV_X1    g0590(.A(new_n751), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G116), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n732), .A2(G87), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n757), .B1(new_n752), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G303), .B2(new_n727), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n742), .A2(new_n797), .B1(new_n722), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n259), .B(new_n799), .C1(G107), .C2(new_n740), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n792), .A2(new_n793), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n719), .A2(G143), .B1(G150), .B2(new_n743), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n803), .B2(new_n726), .C1(new_n751), .C2(new_n760), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT34), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n739), .A2(new_n213), .B1(new_n731), .B2(new_n317), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G132), .B2(new_n723), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n259), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n734), .A2(new_n357), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n801), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n766), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n428), .A2(new_n652), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n422), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n429), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n429), .A2(new_n652), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n768), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n766), .A2(new_n768), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n204), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n811), .A2(new_n775), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n817), .B(KEYINPUT99), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n626), .B2(new_n653), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n652), .B(new_n817), .C1(new_n616), .C2(new_n625), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(new_n702), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n821), .B1(new_n826), .B2(new_n775), .ZN(G384));
  INV_X1    g0627(.A(new_n650), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n365), .A2(new_n367), .ZN(new_n829));
  NOR2_X1   g0629(.A1(KEYINPUT100), .A2(KEYINPUT16), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n387), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n365), .B(new_n367), .C1(KEYINPUT100), .C2(KEYINPUT16), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n351), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n828), .B(new_n834), .C1(new_n635), .C2(new_n638), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n632), .B1(new_n395), .B2(new_n828), .ZN(new_n836));
  INV_X1    g0636(.A(new_n637), .ZN(new_n837));
  XOR2_X1   g0637(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n396), .A2(new_n650), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n637), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n835), .A2(KEYINPUT38), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n839), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n638), .A2(KEYINPUT104), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT104), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n636), .B(new_n849), .C1(new_n347), .C2(new_n637), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n399), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n370), .A2(new_n650), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n844), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n815), .B1(new_n429), .B2(new_n813), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n326), .A2(new_n652), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI221_X4 g0658(.A(new_n858), .B1(new_n332), .B2(new_n333), .C1(new_n316), .C2(new_n326), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n327), .A2(new_n653), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n701), .B2(new_n700), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n835), .A2(KEYINPUT38), .A3(new_n843), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n835), .B2(new_n843), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n327), .A2(new_n334), .A3(new_n857), .ZN(new_n868));
  INV_X1    g0668(.A(new_n860), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n817), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n555), .A2(new_n593), .A3(new_n595), .A4(new_n653), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n695), .A2(new_n698), .A3(new_n652), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n698), .B1(new_n695), .B2(new_n652), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n864), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT107), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n700), .A2(new_n701), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n870), .C1(new_n865), .C2(new_n866), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(KEYINPUT107), .A3(new_n864), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n863), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n432), .A3(new_n879), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n650), .B(new_n833), .C1(new_n392), .C2(new_n399), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n834), .A2(new_n840), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n842), .B1(new_n887), .B2(new_n837), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n845), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n885), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n844), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n877), .B(KEYINPUT40), .C1(new_n891), .C2(new_n862), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT107), .B1(new_n880), .B2(new_n864), .ZN(new_n893));
  OAI211_X1 g0693(.A(G330), .B(new_n884), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n432), .A2(new_n702), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n883), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT108), .Z(new_n898));
  NAND3_X1  g0698(.A1(new_n432), .A2(new_n711), .A3(new_n714), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n643), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(KEYINPUT105), .B(KEYINPUT106), .Z(new_n902));
  XNOR2_X1  g0702(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n859), .A2(new_n860), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n891), .B(new_n905), .C1(new_n824), .C2(new_n815), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n635), .A2(new_n650), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT102), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(KEYINPUT102), .A3(new_n907), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n327), .A2(new_n652), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(new_n844), .C1(new_n853), .C2(new_n854), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n910), .B(new_n911), .C1(new_n913), .C2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n903), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n251), .B2(new_n772), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n536), .B1(new_n438), .B2(KEYINPUT35), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n230), .C1(KEYINPUT35), .C2(new_n438), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT36), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n231), .A2(new_n358), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n924), .A2(new_n216), .B1(G50), .B2(new_n317), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n646), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n920), .A2(new_n923), .A3(new_n926), .ZN(G367));
  AOI22_X1  g0727(.A1(new_n791), .A2(G283), .B1(G317), .B2(new_n723), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n265), .C1(new_n798), .C2(new_n726), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(G107), .B2(new_n735), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n719), .A2(G303), .B1(G294), .B2(new_n743), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n732), .A2(G97), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n740), .A2(G116), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT46), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n751), .A2(new_n213), .B1(new_n760), .B2(new_n742), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n259), .B1(new_n803), .B2(new_n722), .C1(new_n936), .C2(KEYINPUT113), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G58), .B2(new_n740), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n732), .A2(new_n215), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(KEYINPUT113), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n735), .A2(G68), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n752), .B2(new_n283), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n942), .A2(KEYINPUT112), .B1(G143), .B2(new_n727), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT47), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n766), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n509), .A2(new_n517), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n652), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n607), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n622), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n770), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n785), .B1(new_n209), .B2(new_n402), .C1(new_n241), .C2(new_n777), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n948), .A2(new_n775), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n598), .B1(new_n523), .B2(new_n653), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n485), .B2(new_n653), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT110), .Z(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(new_n588), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n652), .B1(new_n964), .B2(new_n485), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n596), .A3(new_n665), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT42), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n958), .B(new_n960), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n965), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n969), .B2(new_n960), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n663), .A2(new_n963), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n970), .B(new_n971), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n773), .A2(G1), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n666), .A2(new_n962), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT45), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n666), .A2(new_n962), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n662), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT111), .ZN(new_n980));
  MUX2_X1   g0780(.A(new_n661), .B(new_n596), .S(new_n665), .Z(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(new_n658), .Z(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(new_n715), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n662), .B2(new_n978), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n715), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n669), .B(KEYINPUT41), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n973), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n957), .B1(new_n972), .B2(new_n987), .ZN(G387));
  INV_X1    g0788(.A(new_n766), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n752), .A2(new_n990), .B1(new_n798), .B2(new_n742), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G322), .B2(new_n727), .ZN(new_n992));
  INV_X1    g0792(.A(G303), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(new_n751), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT48), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n797), .B2(new_n734), .C1(new_n794), .C2(new_n739), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n259), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n723), .A2(G326), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n732), .A2(G116), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT115), .B(G150), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n722), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n738), .A2(G68), .B1(new_n496), .B2(new_n735), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n760), .B2(new_n726), .C1(new_n281), .C2(new_n742), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G50), .C2(new_n719), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n740), .A2(new_n215), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1007), .A2(new_n259), .A3(new_n932), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n989), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G45), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n238), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT114), .Z(new_n1013));
  NOR2_X1   g0813(.A1(new_n281), .A2(G50), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g0815(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n671), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n776), .A3(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(G107), .B2(new_n209), .C1(new_n671), .C2(new_n780), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1019), .A2(new_n785), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n661), .A2(new_n770), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1010), .A2(new_n774), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n982), .B2(new_n973), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n669), .B1(new_n982), .B2(new_n715), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n983), .B2(new_n1024), .ZN(G393));
  XNOR2_X1  g0825(.A(new_n978), .B(new_n663), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n669), .B1(new_n1026), .B2(new_n983), .C1(new_n980), .C2(new_n984), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n785), .B1(new_n222), .B2(new_n209), .C1(new_n249), .C2(new_n777), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n791), .A2(new_n348), .B1(G50), .B2(new_n743), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n734), .A2(new_n204), .ZN(new_n1030));
  INV_X1    g0830(.A(G143), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n259), .B1(new_n722), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G68), .C2(new_n740), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n719), .A2(G159), .B1(new_n727), .B2(G150), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT51), .Z(new_n1035));
  NAND4_X1  g0835(.A1(new_n1029), .A2(new_n793), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n739), .A2(new_n797), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n742), .A2(new_n993), .B1(new_n734), .B2(new_n536), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(G322), .C2(new_n723), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n259), .B1(new_n738), .B2(G294), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n755), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n719), .A2(G311), .B1(new_n727), .B2(G317), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT52), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1036), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT116), .Z(new_n1045));
  OAI211_X1 g0845(.A(new_n775), .B(new_n1028), .C1(new_n1045), .C2(new_n989), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n963), .B2(new_n770), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1026), .B2(new_n973), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1027), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT117), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT117), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1027), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(G390));
  NAND3_X1  g0853(.A1(new_n626), .A2(new_n653), .A3(new_n856), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n904), .B1(new_n1054), .B2(new_n816), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n914), .B(new_n916), .C1(new_n1055), .C2(new_n912), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n855), .A2(new_n913), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n708), .A2(new_n709), .A3(new_n816), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n814), .A3(new_n905), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n702), .A2(new_n870), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1056), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n899), .A2(new_n643), .A3(new_n895), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n702), .A2(new_n856), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1062), .B1(new_n1068), .B2(new_n905), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n815), .B2(new_n824), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1058), .A2(new_n814), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n702), .A2(new_n822), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1062), .C1(new_n905), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1064), .A2(new_n1067), .A3(new_n1065), .A4(new_n1074), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n669), .A3(new_n1077), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1056), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1062), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n973), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n917), .A2(new_n768), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n751), .A2(new_n222), .B1(new_n536), .B2(new_n752), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1084), .A2(new_n1030), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n727), .A2(G283), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n265), .B1(new_n739), .B2(new_n504), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT118), .Z(new_n1088));
  OAI22_X1  g0888(.A1(new_n742), .A2(new_n433), .B1(new_n731), .B2(new_n317), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G294), .B2(new_n723), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  AOI22_X1  g0892(.A1(new_n791), .A2(new_n1092), .B1(G125), .B2(new_n723), .ZN(new_n1093));
  INV_X1    g0893(.A(G128), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n259), .C1(new_n1094), .C2(new_n726), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G159), .B2(new_n735), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n739), .A2(new_n1003), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n719), .A2(G132), .B1(G50), .B2(new_n732), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n742), .A2(new_n803), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1091), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n766), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n819), .A2(new_n281), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1083), .A2(new_n775), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1078), .A2(new_n1082), .A3(new_n1105), .ZN(G378));
  INV_X1    g0906(.A(KEYINPUT57), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n296), .B1(new_n344), .B2(new_n345), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n295), .A2(new_n828), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n296), .B(new_n1109), .C1(new_n344), .C2(new_n345), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1111), .A2(new_n1114), .A3(new_n1112), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n882), .B2(G330), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1118), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n894), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n918), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n911), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT102), .B1(new_n906), .B2(new_n907), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n882), .A2(G330), .A3(new_n1118), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n894), .A2(new_n1120), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n899), .A2(new_n643), .A3(new_n895), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1081), .B2(new_n1074), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1107), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(KEYINPUT57), .A3(new_n1129), .A4(new_n1122), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n669), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1122), .A2(new_n1129), .A3(new_n973), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n774), .B1(new_n1118), .B2(new_n768), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n941), .B1(new_n536), .B2(new_n726), .C1(new_n752), .C2(new_n433), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n259), .B(new_n1139), .C1(new_n496), .C2(new_n738), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n731), .A2(new_n357), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT119), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n467), .A3(new_n1008), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G97), .B2(new_n743), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1140), .B(new_n1144), .C1(new_n797), .C2(new_n722), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT58), .Z(new_n1146));
  OAI21_X1  g0946(.A(new_n213), .B1(new_n263), .B2(G41), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n726), .A2(new_n1148), .B1(new_n734), .B2(new_n283), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n738), .A2(G137), .B1(new_n743), .B2(G132), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1094), .B2(new_n752), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(new_n740), .C2(new_n1092), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1153));
  AOI21_X1  g0953(.A(G33), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n723), .B2(G124), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n760), .C2(new_n731), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1147), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n766), .B1(new_n1146), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n819), .A2(new_n213), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1138), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT121), .B1(new_n1137), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1137), .A2(KEYINPUT121), .A3(new_n1161), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1136), .B1(new_n1162), .B2(new_n1163), .ZN(G375));
  NAND3_X1  g0964(.A1(new_n1131), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1075), .A2(new_n986), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n819), .A2(new_n317), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n905), .B2(new_n769), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n265), .B1(new_n204), .B2(new_n731), .C1(new_n751), .C2(new_n433), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n719), .A2(G283), .B1(new_n496), .B2(new_n735), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n794), .B2(new_n726), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n740), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n993), .B2(new_n722), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1169), .B(new_n1173), .C1(G116), .C2(new_n743), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT122), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n722), .A2(new_n1094), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1142), .B1(new_n213), .B2(new_n734), .C1(new_n283), .C2(new_n748), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n743), .A2(new_n1092), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n752), .B2(new_n803), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n265), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n727), .A2(G132), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n760), .C2(new_n739), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n774), .B(new_n1168), .C1(new_n1183), .C2(new_n766), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1074), .B2(new_n973), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1166), .A2(new_n1185), .ZN(G381));
  NOR2_X1   g0986(.A1(G390), .A2(G387), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(G381), .A2(G384), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1188), .A2(G396), .A3(G393), .A4(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G375), .A2(G378), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(G407));
  NAND2_X1  g0992(.A1(new_n651), .A2(G213), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT123), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1191), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(G213), .ZN(G409));
  OAI211_X1 g0997(.A(new_n1136), .B(G378), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1198));
  INV_X1    g0998(.A(G378), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1137), .A2(new_n1161), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n986), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1130), .A2(new_n1132), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1199), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1195), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT60), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1075), .B(new_n669), .C1(new_n1165), .C2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1165), .A2(new_n1206), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1185), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(G384), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(new_n1194), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1211), .A2(G2897), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT61), .B1(new_n1205), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n1193), .A3(new_n1210), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT124), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1218), .A3(new_n1193), .A4(new_n1210), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT62), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1215), .A2(KEYINPUT62), .A3(new_n1194), .A4(new_n1210), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT126), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1204), .A2(new_n1223), .A3(KEYINPUT62), .A4(new_n1210), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1214), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT127), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(G393), .B(G396), .Z(new_n1229));
  NAND2_X1  g1029(.A1(G390), .A2(G387), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1188), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1188), .B2(new_n1230), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(KEYINPUT127), .B(new_n1214), .C1(new_n1220), .C2(new_n1225), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1228), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1233), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1204), .A2(KEYINPUT63), .A3(new_n1210), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT125), .Z(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT63), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT61), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1215), .A2(new_n1193), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1213), .A2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1236), .A2(new_n1238), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1235), .A2(new_n1243), .ZN(G405));
  XNOR2_X1  g1044(.A(G375), .B(new_n1199), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(new_n1210), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1233), .B(new_n1246), .ZN(G402));
endmodule


