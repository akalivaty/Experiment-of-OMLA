//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(G183gat), .B(G190gat), .C1(KEYINPUT66), .C2(KEYINPUT24), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT65), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT23), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n210), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT25), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n203), .B1(new_n207), .B2(new_n205), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n205), .B2(new_n203), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  OR2_X1    g025(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n227), .A2(KEYINPUT23), .A3(new_n211), .A4(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n221), .A4(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT27), .B(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT28), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G183gat), .ZN(new_n237));
  AND4_X1   g036(.A1(KEYINPUT28), .A2(new_n235), .A3(new_n237), .A4(new_n232), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n203), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n240), .A2(new_n219), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n213), .A2(new_n215), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n217), .B2(new_n242), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n223), .B(new_n230), .C1(new_n239), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G127gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT1), .B1(new_n248), .B2(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(G113gat), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G113gat), .A2(G120gat), .ZN(new_n253));
  INV_X1    g052(.A(G134gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G127gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n249), .A2(new_n252), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(G113gat), .A2(G120gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT70), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n252), .A2(new_n260), .A3(new_n253), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT1), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n254), .B2(G127gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n248), .B2(G134gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n254), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n264), .A2(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n247), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n247), .A2(new_n270), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n247), .B2(new_n270), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n202), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n272), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n247), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n278));
  AND4_X1   g077(.A1(new_n202), .A2(new_n277), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(KEYINPUT33), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT72), .B(new_n285), .C1(new_n274), .C2(new_n275), .ZN(new_n286));
  XOR2_X1   g085(.A(G15gat), .B(G43gat), .Z(new_n287));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT32), .B1(new_n274), .B2(new_n275), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n284), .A2(new_n286), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n289), .A2(KEYINPUT33), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n281), .B1(new_n294), .B2(KEYINPUT73), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n296), .B(new_n280), .C1(new_n291), .C2(new_n293), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT90), .ZN(new_n299));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT31), .B(G50gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G228gat), .A2(G233gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT83), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n307));
  NAND2_X1  g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G204gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G197gat), .ZN(new_n312));
  INV_X1    g111(.A(G197gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G204gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n308), .ZN(new_n316));
  NOR2_X1   g115(.A1(G211gat), .A2(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n307), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n308), .ZN(new_n321));
  XNOR2_X1  g120(.A(G197gat), .B(G204gat), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT84), .A4(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n315), .A2(new_n318), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT2), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n326), .A2(new_n329), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n329), .A2(new_n335), .A3(new_n333), .ZN(new_n336));
  AND2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n334), .B2(new_n340), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n334), .A2(new_n340), .A3(new_n344), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n315), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n320), .A2(new_n353), .A3(new_n308), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n310), .A3(new_n322), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n345), .B1(new_n325), .B2(new_n341), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n343), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n306), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G22gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT3), .B1(new_n356), .B2(new_n349), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n334), .A2(new_n340), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n350), .B2(new_n357), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n356), .B1(new_n349), .B2(new_n348), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n368), .ZN(new_n372));
  INV_X1    g171(.A(new_n304), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n367), .A2(new_n370), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n362), .A2(new_n363), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n363), .B1(new_n362), .B2(new_n374), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n342), .A2(new_n346), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT85), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n371), .B1(new_n360), .B2(new_n343), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n305), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n373), .B1(new_n364), .B2(new_n366), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n350), .A2(new_n368), .A3(new_n357), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n383), .A2(new_n384), .A3(new_n369), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n377), .B(G22gat), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n303), .B1(new_n378), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT88), .ZN(new_n389));
  OAI21_X1  g188(.A(G22gat), .B1(new_n382), .B2(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT87), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n386), .A3(new_n375), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n303), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT89), .B(G22gat), .C1(new_n382), .C2(new_n385), .ZN(new_n396));
  NAND2_X1  g195(.A1(KEYINPUT89), .A2(G22gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n362), .A2(new_n374), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n302), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n299), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  AOI211_X1 g200(.A(KEYINPUT90), .B(new_n401), .C1(new_n389), .C2(new_n394), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n298), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n247), .B2(new_n349), .ZN(new_n406));
  INV_X1    g205(.A(new_n203), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n235), .A2(new_n237), .A3(new_n232), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n231), .A2(KEYINPUT28), .A3(new_n232), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n229), .A2(new_n221), .A3(new_n226), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n225), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n404), .B1(new_n415), .B2(new_n223), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n357), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT75), .B(new_n357), .C1(new_n406), .C2(new_n416), .ZN(new_n420));
  INV_X1    g219(.A(new_n416), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n415), .B2(new_n223), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n421), .B(new_n356), .C1(new_n422), .C2(new_n405), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n419), .A2(new_n420), .A3(new_n423), .A4(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n406), .A2(new_n416), .A3(new_n357), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n418), .B2(new_n417), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n420), .A4(new_n429), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G1gat), .B(G29gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G57gat), .B(G85gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT81), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n439), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n270), .A2(new_n365), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n346), .A2(new_n270), .A3(new_n348), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n448), .C1(KEYINPUT4), .C2(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n450), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n446), .B1(new_n270), .B2(new_n365), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n457), .A2(new_n458), .B1(new_n444), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT77), .B(new_n446), .C1(new_n270), .C2(new_n365), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT79), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n270), .A2(new_n365), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n451), .B1(new_n464), .B2(new_n444), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n453), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n457), .A2(new_n458), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n444), .A2(new_n459), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n461), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n456), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n270), .B(new_n365), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n452), .B1(new_n473), .B2(new_n451), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT79), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n443), .B(new_n455), .C1(new_n467), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n463), .B1(new_n462), .B2(new_n466), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(KEYINPUT79), .A3(new_n474), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n454), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(new_n443), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n481), .A2(new_n477), .A3(new_n443), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n436), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT82), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n455), .B1(new_n467), .B2(new_n475), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n442), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n477), .A3(new_n476), .ZN(new_n489));
  INV_X1    g288(.A(new_n484), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n436), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT35), .B1(new_n403), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n429), .B1(new_n433), .B2(new_n420), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n430), .A2(KEYINPUT30), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n496), .B(new_n435), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n431), .B2(new_n435), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n294), .A2(new_n280), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n281), .A2(new_n291), .A3(new_n293), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n502), .A2(new_n505), .A3(new_n506), .A4(new_n491), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n392), .A2(new_n393), .A3(new_n303), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n393), .B1(new_n392), .B2(new_n303), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n399), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT90), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n395), .A2(new_n299), .A3(new_n399), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n505), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n298), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n400), .A2(new_n402), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n494), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n491), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n424), .A2(KEYINPUT37), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n427), .B1(new_n424), .B2(KEYINPUT37), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT38), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n423), .A2(new_n417), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT38), .B1(new_n524), .B2(KEYINPUT37), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n427), .C1(KEYINPUT37), .C2(new_n424), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n523), .A2(new_n430), .A3(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n511), .A2(new_n512), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT92), .B(KEYINPUT39), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n449), .A2(new_n451), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n449), .A2(new_n451), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT39), .B1(new_n473), .B2(new_n451), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n443), .B(new_n530), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT40), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n531), .B(KEYINPUT39), .C1(new_n451), .C2(new_n473), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n537), .A2(KEYINPUT40), .A3(new_n443), .A4(new_n530), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(new_n482), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n500), .B2(new_n501), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n540), .B(new_n543), .C1(new_n500), .C2(new_n501), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n495), .A2(new_n514), .B1(new_n519), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n549));
  INV_X1    g348(.A(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n552), .A2(new_n553), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n555));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n554), .B2(KEYINPUT15), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT17), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n572), .A3(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n562), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n560), .A2(KEYINPUT17), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n558), .B2(new_n559), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT99), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT95), .Z(new_n585));
  INV_X1    g384(.A(KEYINPUT41), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n576), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n560), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT100), .Z(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(KEYINPUT101), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n577), .B2(new_n582), .ZN(new_n596));
  INV_X1    g395(.A(new_n592), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n586), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT96), .Z(new_n605));
  NAND4_X1  g404(.A1(new_n593), .A2(new_n598), .A3(new_n599), .A4(new_n601), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n603), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G183gat), .B(G211gat), .Z(new_n610));
  XOR2_X1   g409(.A(G57gat), .B(G64gat), .Z(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(G71gat), .A2(G78gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(KEYINPUT94), .A2(KEYINPUT9), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n615), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT16), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(G1gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G15gat), .B(G22gat), .ZN(new_n630));
  MUX2_X1   g429(.A(G1gat), .B(new_n629), .S(new_n630), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G8gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(KEYINPUT21), .B2(new_n619), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n624), .A2(new_n626), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n627), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n627), .B2(new_n636), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n610), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n627), .A2(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n634), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n627), .A2(new_n635), .A3(new_n636), .ZN(new_n642));
  INV_X1    g441(.A(new_n610), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646));
  INV_X1    g445(.A(G230gat), .ZN(new_n647));
  INV_X1    g446(.A(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n619), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n576), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n574), .A2(new_n619), .A3(new_n575), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT102), .Z(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n652), .A2(new_n660), .A3(new_n653), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n653), .A2(new_n660), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n649), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n655), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n659), .B1(new_n655), .B2(new_n664), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n646), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n655), .A2(new_n664), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n658), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G113gat), .B(G141gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT11), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n211), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n313), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT12), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n561), .A2(new_n632), .ZN(new_n678));
  NAND2_X1  g477(.A1(G229gat), .A2(G233gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n633), .A2(new_n560), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n632), .B(new_n560), .Z(new_n685));
  XOR2_X1   g484(.A(new_n679), .B(KEYINPUT13), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n681), .B2(new_n682), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n677), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n678), .A2(new_n680), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(KEYINPUT18), .A3(new_n679), .ZN(new_n691));
  INV_X1    g490(.A(new_n677), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n691), .A2(new_n683), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n672), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n609), .A2(new_n645), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n548), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n491), .A2(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n491), .A2(KEYINPUT104), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n698), .A2(new_n502), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n708), .B2(G8gat), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT16), .B(G8gat), .Z(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n707), .A2(KEYINPUT105), .A3(KEYINPUT42), .A4(new_n710), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n711), .B2(new_n706), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n717), .B(new_n715), .C1(new_n709), .C2(new_n712), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1325gat));
  INV_X1    g520(.A(new_n505), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n698), .A2(G15gat), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n517), .ZN(new_n724));
  OAI21_X1  g523(.A(G15gat), .B1(new_n698), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n511), .A2(new_n512), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n698), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n547), .B2(new_n609), .ZN(new_n732));
  INV_X1    g531(.A(new_n605), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n592), .B(new_n595), .C1(new_n577), .C2(new_n582), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n590), .A2(new_n592), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n594), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n601), .B1(new_n736), .B2(new_n593), .ZN(new_n737));
  INV_X1    g536(.A(new_n606), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n494), .A2(new_n518), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n546), .A2(new_n742), .A3(new_n724), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n486), .A3(new_n493), .A4(new_n298), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n513), .B1(KEYINPUT35), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT44), .B(new_n741), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n732), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n645), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n696), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G29gat), .B1(new_n751), .B2(new_n702), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n547), .A2(new_n609), .A3(new_n749), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n550), .A3(new_n703), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1328gat));
  INV_X1    g555(.A(new_n502), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n551), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT46), .Z(new_n759));
  OAI21_X1  g558(.A(G36gat), .B1(new_n751), .B2(new_n502), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1329gat));
  NAND4_X1  g560(.A1(new_n732), .A2(new_n517), .A3(new_n746), .A4(new_n750), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n722), .A2(G43gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n753), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n763), .A2(KEYINPUT107), .B1(new_n753), .B2(new_n764), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n762), .A2(new_n769), .A3(G43gat), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n767), .B(KEYINPUT47), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n770), .A3(new_n765), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT108), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n766), .B1(new_n771), .B2(new_n775), .ZN(G1330gat));
  OAI21_X1  g575(.A(G50gat), .B1(new_n751), .B2(new_n727), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n727), .A2(G50gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n753), .A2(new_n778), .B1(KEYINPUT109), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n779), .A2(KEYINPUT109), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1331gat));
  NAND4_X1  g582(.A1(new_n739), .A2(new_n645), .A3(new_n740), .A4(new_n695), .ZN(new_n784));
  INV_X1    g583(.A(new_n672), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n548), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n702), .B(KEYINPUT110), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g589(.A(new_n787), .B(KEYINPUT111), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  NOR4_X1   g592(.A1(new_n791), .A2(new_n502), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n791), .A2(new_n502), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n792), .B2(new_n795), .ZN(G1333gat));
  OAI21_X1  g595(.A(G71gat), .B1(new_n791), .B2(new_n724), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n787), .A2(G71gat), .A3(new_n722), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1334gat));
  NOR2_X1   g600(.A1(new_n791), .A2(new_n727), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g602(.A1(new_n785), .A2(new_n645), .A3(new_n694), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n747), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G85gat), .B1(new_n805), .B2(new_n702), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n547), .A2(new_n609), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n645), .A2(new_n694), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT51), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n702), .A2(new_n785), .A3(G85gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT112), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n806), .B(new_n815), .C1(new_n810), .C2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1336gat));
  NAND3_X1  g616(.A1(new_n747), .A2(new_n757), .A3(new_n804), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n785), .A2(G92gat), .A3(new_n502), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n819), .B(new_n820), .C1(new_n810), .C2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT113), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n809), .B(new_n825), .Z(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(new_n821), .B1(G92gat), .B2(new_n818), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n827), .B2(new_n820), .ZN(G1337gat));
  XOR2_X1   g627(.A(KEYINPUT114), .B(G99gat), .Z(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n805), .B2(new_n724), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n785), .A2(new_n722), .A3(new_n829), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n810), .B2(new_n831), .ZN(G1338gat));
  NAND3_X1  g631(.A1(new_n747), .A2(new_n518), .A3(new_n804), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G106gat), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n727), .A2(new_n785), .A3(G106gat), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n834), .B(new_n835), .C1(new_n810), .C2(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n826), .A2(new_n836), .B1(G106gat), .B2(new_n833), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n835), .ZN(G1339gat));
  NOR2_X1   g639(.A1(new_n784), .A2(new_n672), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n659), .B1(new_n663), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n661), .A2(new_n662), .A3(new_n649), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n663), .A3(new_n845), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n664), .A2(KEYINPUT54), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT55), .B(new_n846), .C1(new_n851), .C2(new_n848), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n665), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n676), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n690), .A2(new_n679), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n685), .A2(new_n686), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT115), .A4(new_n665), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n855), .A2(new_n693), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n843), .B1(new_n609), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n741), .A2(new_n863), .A3(KEYINPUT116), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n855), .A2(new_n694), .A3(new_n860), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n693), .A2(new_n859), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n785), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n862), .A2(new_n864), .B1(new_n867), .B2(new_n609), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n842), .B1(new_n868), .B2(new_n645), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n788), .A2(new_n757), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n403), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n694), .ZN(new_n874));
  INV_X1    g673(.A(new_n869), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n703), .A2(new_n502), .A3(new_n505), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n518), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n695), .A2(new_n250), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1340gat));
  AOI21_X1  g678(.A(G120gat), .B1(new_n873), .B2(new_n672), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n785), .A2(new_n251), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n877), .B2(new_n881), .ZN(G1341gat));
  NAND3_X1  g681(.A1(new_n873), .A2(new_n248), .A3(new_n645), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n877), .A2(new_n645), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n248), .B2(new_n884), .ZN(G1342gat));
  NAND2_X1  g684(.A1(new_n871), .A2(new_n741), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(G134gat), .A3(new_n403), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n877), .A2(new_n741), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G134gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1343gat));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n702), .A2(new_n757), .A3(new_n517), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT117), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n695), .A2(new_n327), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n869), .B2(new_n518), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n518), .A2(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n862), .A2(new_n864), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n853), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT118), .A4(new_n665), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n695), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n866), .B1(new_n668), .B2(new_n671), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n740), .B(new_n739), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n748), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n897), .B1(new_n906), .B2(new_n842), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n517), .A2(new_n727), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n869), .A2(new_n694), .A3(new_n870), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n327), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n892), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT119), .B(KEYINPUT58), .C1(new_n908), .C2(new_n911), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n914), .A2(new_n915), .B1(new_n913), .B2(new_n912), .ZN(G1344gat));
  XNOR2_X1  g715(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n894), .A2(new_n672), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n853), .A2(new_n866), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n607), .B2(new_n608), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n900), .A2(new_n901), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n903), .B1(new_n923), .B2(new_n694), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n924), .B2(new_n741), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n841), .B1(new_n925), .B2(new_n748), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n919), .B(new_n920), .C1(new_n926), .C2(new_n727), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n645), .B1(new_n904), .B2(new_n922), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n518), .B1(new_n929), .B2(new_n841), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n919), .B1(new_n930), .B2(new_n920), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n867), .A2(new_n609), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n645), .B1(new_n898), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT57), .B(new_n518), .C1(new_n934), .C2(new_n841), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n918), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(KEYINPUT122), .B(new_n917), .C1(new_n936), .C2(new_n328), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n930), .A2(new_n920), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT121), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n935), .A3(new_n927), .ZN(new_n941));
  INV_X1    g740(.A(new_n918), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n328), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n917), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n328), .A2(KEYINPUT59), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n894), .B1(new_n896), .B2(new_n907), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(new_n785), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n937), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n871), .A2(new_n328), .A3(new_n672), .A4(new_n909), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1345gat));
  OAI21_X1  g750(.A(G155gat), .B1(new_n947), .B2(new_n748), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n871), .A2(new_n330), .A3(new_n645), .A4(new_n909), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1346gat));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n947), .B2(new_n609), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G162gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n947), .A2(new_n955), .A3(new_n609), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n909), .A2(new_n331), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n957), .A2(new_n958), .B1(new_n886), .B2(new_n959), .ZN(G1347gat));
  AND2_X1   g759(.A1(new_n788), .A2(new_n757), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n869), .A2(new_n961), .A3(new_n727), .A4(new_n505), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n211), .A3(new_n695), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n872), .A2(new_n757), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n875), .A2(new_n703), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n694), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n963), .B1(new_n966), .B2(new_n211), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n965), .B2(new_n672), .ZN(new_n968));
  INV_X1    g767(.A(new_n962), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n785), .B1(new_n227), .B2(new_n228), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(G1349gat));
  NAND3_X1  g770(.A1(new_n965), .A2(new_n231), .A3(new_n645), .ZN(new_n972));
  OAI21_X1  g771(.A(G183gat), .B1(new_n962), .B2(new_n748), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n965), .A2(new_n232), .A3(new_n741), .ZN(new_n976));
  OAI21_X1  g775(.A(G190gat), .B1(new_n962), .B2(new_n609), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n977), .A2(KEYINPUT61), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n977), .A2(KEYINPUT61), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1351gat));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n724), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n941), .A2(new_n694), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(KEYINPUT125), .B(G197gat), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n875), .A2(new_n703), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n909), .A2(new_n757), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT124), .Z(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n694), .A2(new_n984), .ZN(new_n989));
  OAI22_X1  g788(.A1(new_n983), .A2(new_n984), .B1(new_n988), .B2(new_n989), .ZN(G1352gat));
  NAND3_X1  g789(.A1(new_n941), .A2(new_n672), .A3(new_n982), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n311), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(new_n992), .B2(new_n991), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n985), .A2(new_n311), .A3(new_n672), .A4(new_n987), .ZN(new_n995));
  XOR2_X1   g794(.A(new_n995), .B(KEYINPUT62), .Z(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1353gat));
  OR3_X1    g796(.A1(new_n988), .A2(G211gat), .A3(new_n748), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n941), .A2(new_n645), .A3(new_n982), .ZN(new_n999));
  AND3_X1   g798(.A1(new_n999), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT63), .B1(new_n999), .B2(G211gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G1354gat));
  NAND3_X1  g801(.A1(new_n941), .A2(new_n741), .A3(new_n982), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G218gat), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n609), .A2(G218gat), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n985), .A2(new_n987), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT127), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1004), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1010), .ZN(G1355gat));
endmodule


