//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT66), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n480), .A2(new_n482), .A3(new_n475), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n475), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n495), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n481), .A2(G126), .A3(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n481), .B2(new_n505), .ZN(new_n506));
  AND4_X1   g081(.A1(new_n503), .A2(new_n505), .A3(new_n465), .A4(new_n467), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n501), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(new_n514), .B1(new_n511), .B2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n511), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n519), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n518), .A2(G51), .ZN(new_n529));
  AND3_X1   g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n515), .A2(new_n516), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT69), .B(G89), .Z(new_n532));
  OAI221_X1 g107(.A(new_n529), .B1(KEYINPUT7), .B2(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(G63), .ZN(new_n535));
  NAND3_X1  g110(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n534), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n516), .A2(G543), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n531), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n534), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n531), .A2(new_n548), .B1(new_n549), .B2(new_n543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n516), .A2(KEYINPUT70), .A3(G53), .A4(G543), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n558), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT71), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g141(.A(KEYINPUT72), .B(G65), .Z(new_n567));
  AOI22_X1  g142(.A1(new_n515), .A2(new_n567), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n534), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n560), .A2(KEYINPUT71), .A3(KEYINPUT9), .A4(new_n561), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n517), .A2(G91), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(G299));
  OR2_X1    g147(.A1(new_n540), .A2(new_n544), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  OAI21_X1  g149(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n518), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n515), .A2(G87), .A3(new_n516), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT73), .Z(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n534), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n531), .A2(new_n583), .B1(new_n584), .B2(new_n543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n517), .A2(G85), .B1(G47), .B2(new_n518), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n523), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n515), .A2(G92), .A3(new_n516), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n523), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n594), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n594), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G299), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(G168), .ZN(G280));
  XOR2_X1   g183(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n484), .A2(G123), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT76), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n464), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n487), .A2(G135), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G14), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT78), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT17), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n646), .B2(new_n648), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n648), .A3(new_n651), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2100), .Z(G227));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n669), .C2(new_n668), .ZN(new_n672));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT79), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  OR2_X1    g256(.A1(G95), .A2(G2105), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n682), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n683));
  INV_X1    g258(.A(G119), .ZN(new_n684));
  INV_X1    g259(.A(G131), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n683), .B1(new_n483), .B2(new_n684), .C1(new_n685), .C2(new_n486), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(KEYINPUT80), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(KEYINPUT80), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(G25), .B(new_n689), .S(G29), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT35), .B(G1991), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT81), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G24), .B(G290), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT82), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  AND2_X1   g271(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G22), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G166), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT85), .B(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(G16), .B2(G23), .ZN(new_n703));
  OR3_X1    g278(.A1(KEYINPUT83), .A2(G16), .A3(G23), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n704), .C1(new_n578), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT84), .B(KEYINPUT33), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(G6), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n586), .B2(new_n705), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n702), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT34), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n698), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n698), .B(new_n715), .C1(KEYINPUT86), .C2(KEYINPUT36), .ZN(new_n719));
  NAND2_X1  g294(.A1(G299), .A2(G16), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G20), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1956), .Z(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2090), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT94), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G34), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n477), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G164), .A2(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G27), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT92), .B(G28), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT30), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n743), .A2(new_n744), .B1(new_n727), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(G29), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n484), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n487), .A2(G141), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND4_X1  g328(.A1(new_n749), .A2(new_n750), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n727), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G5), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G171), .B2(G16), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n741), .B(new_n758), .C1(G1961), .C2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n730), .A2(G2090), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n743), .A2(new_n744), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT31), .B(G11), .Z(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G4), .B2(G16), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n766), .A2(G4), .A3(G16), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n602), .C2(new_n705), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1348), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n761), .A2(new_n762), .A3(new_n765), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G21), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G168), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT91), .B(G1966), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n727), .B2(new_n623), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n727), .A2(G26), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n779));
  INV_X1    g354(.A(G140), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n486), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G128), .B2(new_n484), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n777), .B1(new_n782), .B2(new_n727), .ZN(new_n783));
  MUX2_X1   g358(.A(new_n777), .B(new_n783), .S(KEYINPUT28), .Z(new_n784));
  INV_X1    g359(.A(G2072), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n727), .A2(G33), .ZN(new_n786));
  NAND2_X1  g361(.A1(G115), .A2(G2104), .ZN(new_n787));
  INV_X1    g362(.A(G127), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n468), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2105), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT25), .Z(new_n792));
  INV_X1    g367(.A(G139), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n792), .C1(new_n486), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT89), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n786), .B1(new_n795), .B2(G29), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n784), .A2(G2067), .B1(new_n785), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G2067), .B2(new_n784), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n771), .A2(new_n776), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n718), .A2(new_n719), .A3(new_n733), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n739), .A2(new_n740), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n801), .B1(new_n760), .B2(G1961), .C1(new_n755), .C2(new_n756), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT93), .Z(new_n803));
  NOR2_X1   g378(.A1(new_n796), .A2(new_n785), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT90), .Z(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G19), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n551), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT88), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1341), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n800), .A2(new_n803), .A3(new_n805), .A4(new_n810), .ZN(G311));
  INV_X1    g386(.A(new_n800), .ZN(new_n812));
  INV_X1    g387(.A(new_n803), .ZN(new_n813));
  INV_X1    g388(.A(new_n805), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n809), .ZN(G150));
  AOI22_X1  g390(.A1(new_n517), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n523), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G651), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n603), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT39), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n547), .A2(new_n550), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n826), .A2(KEYINPUT96), .A3(new_n821), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n816), .A2(new_n828), .A3(new_n820), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n531), .A2(new_n830), .B1(new_n831), .B2(new_n543), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n515), .A2(G67), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n534), .B1(new_n833), .B2(new_n817), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT96), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n829), .A2(new_n835), .A3(new_n551), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n825), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n823), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT97), .ZN(G145));
  INV_X1    g418(.A(new_n623), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n689), .B(new_n754), .Z(new_n845));
  OR2_X1    g420(.A1(G106), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n847));
  INV_X1    g422(.A(G130), .ZN(new_n848));
  INV_X1    g423(.A(G142), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n847), .B1(new_n483), .B2(new_n848), .C1(new_n849), .C2(new_n486), .ZN(new_n850));
  INV_X1    g425(.A(new_n626), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n484), .A2(G130), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n487), .A2(G142), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n626), .A4(new_n847), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G164), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n852), .A2(new_n508), .A3(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n782), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n795), .A2(KEYINPUT98), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n795), .B2(KEYINPUT98), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n865), .A2(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n845), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n859), .B1(new_n863), .B2(new_n862), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n689), .B(new_n754), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n865), .A2(new_n861), .A3(new_n858), .A4(new_n857), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n491), .B(new_n477), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n867), .A2(new_n872), .A3(new_n868), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n844), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT99), .B(G37), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n844), .A3(new_n877), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n821), .A2(new_n606), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n837), .B(new_n612), .ZN(new_n886));
  OR2_X1    g461(.A1(G299), .A2(new_n602), .ZN(new_n887));
  NAND2_X1  g462(.A1(G299), .A2(new_n602), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(new_n888), .ZN(new_n892));
  NOR2_X1   g467(.A1(G299), .A2(new_n602), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(KEYINPUT41), .A3(new_n888), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n890), .B1(new_n886), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  XNOR2_X1  g473(.A(G290), .B(KEYINPUT101), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n519), .A2(new_n578), .A3(new_n526), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n578), .B1(new_n519), .B2(new_n526), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n586), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n578), .ZN(new_n904));
  NAND2_X1  g479(.A1(G303), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G305), .B1(new_n905), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n899), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  XNOR2_X1  g483(.A(G290), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n586), .B1(new_n901), .B2(new_n902), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(G305), .A3(new_n900), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n898), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n885), .B1(new_n914), .B2(new_n606), .ZN(G295));
  OAI21_X1  g490(.A(new_n885), .B1(new_n914), .B2(new_n606), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND2_X1  g492(.A1(G168), .A2(G301), .ZN(new_n918));
  OAI21_X1  g493(.A(G171), .B1(new_n537), .B2(new_n533), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n837), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n918), .A2(new_n827), .A3(new_n836), .A4(new_n919), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n894), .A2(new_n895), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n892), .A2(new_n893), .ZN(new_n924));
  AND4_X1   g499(.A1(new_n827), .A2(new_n918), .A3(new_n836), .A4(new_n919), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n918), .A2(new_n919), .B1(new_n827), .B2(new_n836), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n917), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n922), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT104), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n913), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n913), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n907), .A2(new_n912), .A3(KEYINPUT105), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n923), .A2(new_n927), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n932), .A2(new_n881), .A3(new_n934), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n928), .B2(new_n930), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n942), .A2(KEYINPUT106), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT106), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n931), .A2(new_n913), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(new_n947), .B2(new_n934), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n944), .A2(new_n945), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n934), .A4(new_n932), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n943), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n942), .A2(KEYINPUT106), .A3(new_n943), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n934), .A3(new_n932), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n932), .A2(new_n940), .A3(new_n881), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G2067), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n782), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n689), .A2(new_n691), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n754), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n860), .A2(G2067), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n966), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n508), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(KEYINPUT108), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(KEYINPUT108), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT45), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n974), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n974), .ZN(new_n982));
  OR2_X1    g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n985));
  XNOR2_X1  g560(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n689), .A2(new_n691), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n972), .A2(new_n987), .A3(new_n967), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n982), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n981), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n980), .A2(new_n969), .A3(new_n974), .ZN(new_n991));
  NAND2_X1  g566(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n971), .A2(new_n966), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(new_n754), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n982), .A2(new_n995), .B1(KEYINPUT124), .B2(KEYINPUT46), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT125), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(KEYINPUT47), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n990), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT113), .B(G1981), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n586), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n586), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT114), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(KEYINPUT114), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1006), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n579), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(new_n1004), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n976), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G166), .A2(new_n1018), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n1024));
  OAI22_X1  g599(.A1(G166), .A2(new_n1018), .B1(KEYINPUT112), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n508), .A2(KEYINPUT50), .A3(new_n975), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT50), .B1(new_n508), .B2(new_n975), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n974), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(KEYINPUT111), .A3(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n501), .A2(new_n502), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n506), .A2(new_n507), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT45), .B(new_n975), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT109), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n976), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n1041), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n974), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1043), .A2(KEYINPUT110), .A3(new_n974), .A4(new_n1044), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(G8), .B(new_n1026), .C1(new_n1036), .C2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1011), .B(new_n1019), .C1(new_n1006), .C2(new_n1010), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n578), .A2(new_n1013), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1020), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT52), .B1(new_n1020), .B2(new_n1053), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1015), .A2(new_n1020), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1032), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1026), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n740), .B(new_n974), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n508), .B2(new_n975), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1016), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1064), .B1(new_n1067), .B2(G1966), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1068), .B2(G286), .ZN(new_n1069));
  OAI211_X1 g644(.A(G168), .B(new_n1064), .C1(new_n1067), .C2(G1966), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1063), .B1(new_n1070), .B2(G8), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT62), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1057), .ZN(new_n1075));
  AND4_X1   g650(.A1(new_n1062), .A2(new_n1074), .A3(new_n1050), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1073), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1071), .B2(new_n1069), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(KEYINPUT62), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1047), .A2(new_n744), .A3(new_n1048), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1030), .A2(G1961), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1067), .A2(KEYINPUT53), .A3(new_n744), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G171), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1079), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1058), .B1(new_n1076), .B2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1068), .A2(G8), .A3(G168), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1062), .A2(new_n1050), .A3(new_n1075), .A4(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1036), .B2(new_n1049), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1061), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(new_n1050), .A3(new_n1075), .A4(new_n1091), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1090), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1062), .A2(new_n1050), .A3(new_n1075), .A4(new_n1078), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1030), .A2(G1961), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1016), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1039), .C1(KEYINPUT122), .C2(G2078), .ZN(new_n1105));
  OR3_X1    g680(.A1(new_n980), .A2(new_n1081), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(G301), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT54), .B1(new_n1088), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1082), .A2(G301), .A3(new_n1086), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(KEYINPUT123), .A3(KEYINPUT54), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(KEYINPUT54), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1101), .B(new_n1108), .C1(new_n1112), .C2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1043), .A2(new_n974), .A3(new_n1044), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT116), .B(G1956), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1029), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G299), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1122), .B2(new_n1120), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(KEYINPUT61), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1123), .A2(new_n1130), .A3(new_n1126), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1118), .A2(new_n969), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n976), .B2(new_n1016), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n826), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT59), .Z(new_n1137));
  NAND3_X1  g712(.A1(new_n1017), .A2(KEYINPUT118), .A3(new_n965), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n974), .A2(new_n975), .A3(new_n965), .A4(new_n508), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G1348), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1029), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1144), .A3(KEYINPUT119), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n603), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1148), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT119), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT60), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(KEYINPUT121), .A3(new_n602), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1154), .A2(new_n1158), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1132), .B(new_n1137), .C1(new_n1150), .C2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1123), .B(KEYINPUT120), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n1126), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1149), .A2(new_n602), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1127), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1100), .B1(new_n1117), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n988), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(G1986), .B2(G290), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n982), .B1(new_n1168), .B2(new_n983), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1002), .B1(new_n1166), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(new_n941), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n956), .A2(new_n932), .A3(new_n957), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1173), .B2(new_n933), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n875), .A2(new_n844), .A3(new_n877), .ZN(new_n1175));
  NOR3_X1   g749(.A1(new_n1175), .A2(new_n878), .A3(new_n880), .ZN(new_n1176));
  NOR2_X1   g750(.A1(G227), .A2(new_n461), .ZN(new_n1177));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n1178));
  OAI21_X1  g752(.A(new_n643), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n1180), .A2(new_n680), .A3(new_n679), .ZN(new_n1181));
  NOR4_X1   g755(.A1(new_n1174), .A2(new_n1176), .A3(new_n1179), .A4(new_n1181), .ZN(G308));
  INV_X1    g756(.A(new_n1179), .ZN(new_n1183));
  INV_X1    g757(.A(new_n1181), .ZN(new_n1184));
  NAND4_X1  g758(.A1(new_n948), .A2(new_n883), .A3(new_n1183), .A4(new_n1184), .ZN(G225));
endmodule


