//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n193), .A2(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n191), .A2(G143), .ZN(new_n203));
  OAI211_X1 g017(.A(G128), .B(new_n201), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n192), .B(new_n194), .C1(KEYINPUT1), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n200), .B1(new_n208), .B2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G224), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G953), .ZN(new_n211));
  XOR2_X1   g025(.A(new_n209), .B(new_n211), .Z(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G116), .ZN(new_n214));
  OAI21_X1  g028(.A(G113), .B1(new_n214), .B2(KEYINPUT5), .ZN(new_n215));
  XNOR2_X1  g029(.A(G116), .B(G119), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(KEYINPUT5), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G113), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT74), .B(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n224), .B2(G107), .ZN(new_n225));
  AOI21_X1  g039(.A(G101), .B1(new_n224), .B2(G107), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT75), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n225), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(KEYINPUT74), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT74), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G104), .ZN(new_n238));
  AOI21_X1  g052(.A(G107), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(G104), .B1(new_n230), .B2(new_n232), .ZN(new_n240));
  OAI21_X1  g054(.A(G101), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n234), .A2(new_n235), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n235), .B1(new_n234), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n223), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT80), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n238), .A3(G107), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n233), .B(new_n247), .C1(new_n239), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n237), .A2(G104), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n227), .A2(KEYINPUT74), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n229), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT75), .B(G107), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n255), .A2(KEYINPUT3), .B1(new_n256), .B2(new_n228), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n257), .A2(new_n226), .B1(new_n249), .B2(G101), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n252), .B1(new_n258), .B2(new_n246), .ZN(new_n259));
  INV_X1    g073(.A(G116), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G119), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n214), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n221), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n233), .B1(new_n239), .B2(new_n248), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n247), .A2(new_n251), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n241), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT76), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n234), .A2(new_n235), .A3(new_n241), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n223), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G122), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n245), .A2(new_n266), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT6), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n245), .A2(new_n266), .A3(new_n274), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n280), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n212), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n275), .B(KEYINPUT8), .Z(new_n286));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n215), .A2(new_n287), .B1(new_n216), .B2(KEYINPUT5), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n287), .B2(new_n215), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n272), .A2(new_n221), .A3(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n290), .A2(KEYINPUT83), .ZN(new_n291));
  OAI22_X1  g105(.A1(G104), .A2(new_n256), .B1(new_n224), .B2(G107), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n257), .A2(new_n226), .B1(G101), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(new_n223), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n290), .B2(KEYINPUT83), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n286), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT7), .B1(new_n210), .B2(G953), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n209), .B(new_n297), .Z(new_n298));
  NAND2_X1  g112(.A1(new_n276), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n285), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n190), .B1(new_n284), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n212), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n276), .A2(KEYINPUT6), .B1(new_n278), .B2(new_n280), .ZN(new_n303));
  INV_X1    g117(.A(new_n283), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n295), .ZN(new_n306));
  INV_X1    g120(.A(new_n286), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n299), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n310), .A3(new_n189), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G214), .B1(G237), .B2(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G237), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G214), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n193), .ZN(new_n318));
  NOR2_X1   g132(.A1(G237), .A2(G953), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT18), .A3(G131), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(new_n191), .ZN(new_n324));
  NAND2_X1  g138(.A1(KEYINPUT18), .A2(G131), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n323), .B2(KEYINPUT16), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n318), .B2(new_n320), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(G146), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n318), .A2(new_n333), .A3(new_n320), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n338), .A2(new_n334), .A3(KEYINPUT17), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n327), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G113), .B(G122), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n227), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n342), .A2(KEYINPUT87), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n343), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n285), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G475), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n336), .B1(new_n338), .B2(new_n334), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n323), .A2(KEYINPUT85), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT19), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n323), .A2(KEYINPUT85), .A3(KEYINPUT19), .ZN(new_n352));
  AOI21_X1  g166(.A(G146), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n327), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n342), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT86), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n342), .B(new_n327), .C1(new_n337), .C2(new_n339), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n354), .A2(KEYINPUT86), .A3(new_n355), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  NOR2_X1   g176(.A1(G475), .A2(G902), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n361), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n347), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G952), .A3(new_n316), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT89), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT21), .B(G898), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(G902), .A3(G953), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT13), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n205), .B2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n205), .A2(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n193), .A2(G128), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n377), .ZN(new_n382));
  OAI21_X1  g196(.A(G134), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G134), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G116), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n260), .A2(G122), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(new_n256), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n256), .A2(new_n387), .A3(new_n388), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n383), .B(new_n385), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n379), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G134), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n385), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n260), .A2(KEYINPUT14), .A3(G122), .ZN(new_n397));
  OAI211_X1 g211(.A(G107), .B(new_n397), .C1(new_n389), .C2(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(new_n256), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT9), .B(G234), .ZN(new_n402));
  INV_X1    g216(.A(G217), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n402), .A2(new_n403), .A3(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT88), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n401), .A2(new_n405), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n285), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n410), .A2(KEYINPUT15), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n376), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n314), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G221), .B1(new_n402), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G469), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT11), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n384), .B2(G137), .ZN(new_n419));
  INV_X1    g233(.A(G137), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT11), .A3(G134), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n384), .A2(G137), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G131), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(new_n421), .A3(new_n333), .A4(new_n422), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n242), .A2(new_n243), .A3(new_n208), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n269), .A2(new_n207), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n430), .A2(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(KEYINPUT78), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT10), .B1(new_n293), .B2(new_n208), .ZN(new_n434));
  INV_X1    g248(.A(new_n199), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n259), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n426), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n208), .A2(KEYINPUT10), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT77), .B1(new_n272), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n441), .B(new_n438), .C1(new_n270), .C2(new_n271), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n436), .B(new_n437), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n428), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n272), .B2(new_n208), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(KEYINPUT78), .A3(new_n430), .A4(new_n426), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT73), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n316), .A2(G227), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n433), .A2(new_n443), .A3(new_n446), .A4(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n436), .B1(new_n440), .B2(new_n442), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n426), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n455), .B2(new_n443), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n417), .B(new_n285), .C1(new_n453), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n443), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n439), .B1(new_n242), .B2(new_n243), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n441), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n272), .A2(KEYINPUT77), .A3(new_n439), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n437), .B1(new_n464), .B2(new_n436), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n450), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n452), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(KEYINPUT79), .A3(new_n417), .A4(new_n285), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n433), .A2(new_n443), .A3(new_n446), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n450), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n455), .A2(new_n443), .A3(new_n451), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n417), .B1(new_n473), .B2(new_n285), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n416), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n319), .A2(G210), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT27), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT26), .B(G101), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n478), .B(KEYINPUT27), .ZN(new_n483));
  INV_X1    g297(.A(new_n481), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n426), .A2(new_n435), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT64), .B1(new_n384), .B2(G137), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT64), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n420), .A3(G134), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n490), .A3(new_n422), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G131), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n425), .A3(new_n206), .A4(new_n204), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n221), .A2(KEYINPUT65), .A3(new_n264), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT65), .B1(new_n221), .B2(new_n264), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n487), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n204), .A2(new_n425), .A3(new_n206), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n491), .A2(G131), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n199), .B1(new_n425), .B2(new_n424), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n265), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n501), .A3(KEYINPUT67), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  INV_X1    g317(.A(new_n265), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n487), .B2(new_n493), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n204), .A2(new_n425), .A3(new_n206), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n509), .A2(new_n492), .B1(new_n426), .B2(new_n435), .ZN(new_n510));
  INV_X1    g324(.A(new_n495), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n221), .A2(new_n264), .A3(KEYINPUT65), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n486), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT30), .B1(new_n499), .B2(new_n500), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n487), .A2(new_n518), .A3(new_n493), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n482), .A2(new_n485), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n510), .B2(new_n513), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n265), .A2(new_n520), .B1(new_n522), .B2(KEYINPUT66), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n487), .A2(new_n493), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n494), .A2(new_n495), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n486), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(KEYINPUT31), .A3(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT30), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n518), .B1(new_n487), .B2(new_n493), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n265), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n496), .A2(KEYINPUT66), .A3(new_n486), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n516), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n477), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n508), .A2(new_n515), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n521), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT31), .B1(new_n523), .B2(new_n528), .ZN(new_n543));
  AND4_X1   g357(.A1(KEYINPUT31), .A2(new_n528), .A3(new_n532), .A4(new_n533), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT32), .A3(new_n538), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n524), .A2(new_n525), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n496), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n514), .B1(new_n548), .B2(KEYINPUT28), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n521), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n520), .A2(new_n265), .B1(new_n510), .B2(new_n513), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n550), .B1(new_n553), .B2(new_n486), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n521), .B(new_n514), .C1(new_n502), .C2(new_n507), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G472), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n540), .A2(new_n546), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n403), .B1(G234), .B2(new_n285), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n205), .A2(G119), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n561), .B1(KEYINPUT72), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n213), .A2(G128), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT72), .B(KEYINPUT23), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n561), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G110), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n330), .A2(G146), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n331), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n561), .A2(KEYINPUT69), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n205), .A3(G119), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n564), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n570), .A2(KEYINPUT70), .A3(new_n564), .A4(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT24), .B(G110), .Z(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT71), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT71), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n575), .A2(new_n581), .A3(new_n576), .A4(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n569), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n323), .A2(new_n191), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n336), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n577), .A2(new_n579), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n566), .A2(G110), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n316), .A2(G221), .A3(G234), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n590), .B(new_n591), .Z(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n592), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n583), .B2(new_n588), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n285), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT25), .A4(new_n285), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n560), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n593), .A2(new_n595), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(G902), .A3(new_n559), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n558), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n414), .A2(new_n476), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n545), .A2(new_n538), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n537), .B2(G902), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT90), .B1(new_n476), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n474), .B1(new_n459), .B2(new_n468), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT90), .ZN(new_n614));
  NOR4_X1   g428(.A1(new_n613), .A2(new_n614), .A3(new_n416), .A4(new_n610), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n313), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT91), .B1(new_n305), .B2(new_n310), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n187), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n284), .B2(new_n300), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n305), .A2(new_n310), .A3(KEYINPUT91), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n188), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT92), .B1(new_n401), .B2(new_n405), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n407), .A2(new_n408), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n401), .A2(new_n405), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT92), .A3(KEYINPUT33), .A4(new_n406), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n627), .A2(new_n629), .A3(G478), .A4(new_n285), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT93), .B(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n409), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n367), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n375), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n624), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n375), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n365), .A2(KEYINPUT94), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n361), .A2(new_n363), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT20), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n364), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n646), .B2(KEYINPUT94), .ZN(new_n647));
  INV_X1    g461(.A(new_n347), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(new_n412), .A3(new_n648), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n642), .A2(new_n619), .A3(new_n623), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n616), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G107), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n609), .A2(new_n608), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n600), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n594), .A2(KEYINPUT36), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n589), .B(new_n658), .Z(new_n659));
  NOR2_X1   g473(.A1(new_n559), .A2(G902), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(KEYINPUT96), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n663));
  INV_X1    g477(.A(new_n661), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n600), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n414), .A2(new_n476), .A3(new_n656), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n371), .B1(new_n670), .B2(new_n374), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n619), .A2(new_n623), .A3(new_n649), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT97), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n666), .A2(new_n558), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n613), .A3(new_n416), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XNOR2_X1  g494(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n671), .B(new_n681), .Z(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n476), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n312), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n301), .A2(KEYINPUT38), .A3(new_n311), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n534), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n521), .B2(new_n548), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n540), .A2(new_n546), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n412), .B1(new_n646), .B2(new_n347), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n666), .A2(new_n617), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n691), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n685), .A2(new_n686), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n193), .ZN(G45));
  INV_X1    g515(.A(new_n624), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT99), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n633), .B1(new_n646), .B2(new_n347), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n703), .B1(new_n704), .B2(new_n672), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n703), .A2(new_n367), .A3(new_n634), .A4(new_n672), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n702), .A2(KEYINPUT100), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT100), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n705), .A2(new_n706), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n709), .B1(new_n624), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n711), .A3(new_n678), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n466), .B2(new_n452), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(new_n417), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n285), .B1(new_n453), .B2(new_n456), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT101), .A3(G469), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n469), .A3(new_n415), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(new_n469), .A3(KEYINPUT102), .A4(new_n415), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n638), .A3(new_n605), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n650), .A3(new_n605), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR2_X1   g542(.A1(new_n677), .A2(new_n413), .ZN(new_n729));
  INV_X1    g543(.A(new_n720), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n702), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NOR2_X1   g546(.A1(new_n624), .A2(new_n697), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n543), .A2(new_n544), .B1(new_n486), .B2(new_n549), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n538), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n609), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n603), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n375), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n722), .A2(new_n733), .A3(new_n723), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NAND2_X1  g554(.A1(new_n666), .A2(new_n736), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n730), .A2(new_n702), .A3(new_n707), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(new_n603), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n546), .A2(new_n557), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT32), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n608), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n301), .A2(new_n311), .A3(new_n313), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n476), .A2(new_n707), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n613), .A2(new_n750), .A3(new_n604), .A4(new_n416), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n752), .A2(KEYINPUT42), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NOR3_X1   g570(.A1(new_n613), .A2(new_n416), .A3(new_n750), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n605), .A3(new_n649), .A4(new_n672), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  INV_X1    g574(.A(new_n473), .ZN(new_n761));
  OAI21_X1  g575(.A(G469), .B1(new_n761), .B2(KEYINPUT45), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n471), .A2(KEYINPUT45), .A3(new_n472), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n417), .A2(new_n285), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n469), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n764), .A2(new_n760), .A3(new_n765), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n415), .A3(new_n683), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n750), .B(KEYINPUT104), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n634), .A2(new_n646), .A3(new_n347), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n775), .B2(KEYINPUT103), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n777), .A3(KEYINPUT43), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n666), .A2(new_n776), .A3(new_n655), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  OR4_X1    g596(.A1(new_n771), .A2(new_n772), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n766), .A2(new_n469), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n415), .B1(new_n785), .B2(new_n768), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(KEYINPUT105), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(KEYINPUT105), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n789), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n770), .A2(new_n415), .A3(new_n791), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n710), .A2(new_n558), .A3(new_n603), .A4(new_n750), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NOR4_X1   g609(.A1(new_n745), .A2(new_n416), .A3(new_n774), .A4(new_n617), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n719), .A2(new_n469), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT106), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n695), .B(new_n691), .C1(new_n798), .C2(new_n797), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n664), .A2(new_n600), .A3(new_n671), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n733), .A2(new_n476), .A3(new_n695), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n679), .A2(new_n712), .A3(new_n743), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT52), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n807));
  INV_X1    g621(.A(new_n412), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n376), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n314), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n612), .A2(new_n615), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n667), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT107), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n457), .A2(new_n458), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT79), .B1(new_n715), .B2(new_n417), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n475), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n415), .A3(new_n611), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n614), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n476), .A2(KEYINPUT90), .A3(new_n611), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n810), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n667), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n314), .A2(new_n637), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n814), .A2(new_n606), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n724), .A2(new_n739), .A3(new_n731), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n817), .A2(new_n415), .A3(new_n707), .A4(new_n751), .ZN(new_n828));
  INV_X1    g642(.A(new_n749), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT42), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n753), .A2(new_n754), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n830), .A2(new_n831), .A3(new_n758), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT108), .B1(new_n828), .B2(new_n741), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n757), .A2(new_n834), .A3(new_n707), .A4(new_n742), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n412), .A2(new_n347), .A3(new_n672), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n677), .A2(new_n647), .A3(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n833), .A2(new_n835), .B1(new_n757), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n827), .A2(new_n832), .A3(new_n727), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n807), .B1(new_n826), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n757), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n755), .A3(new_n758), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n724), .A2(new_n739), .A3(new_n727), .A4(new_n731), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n822), .B1(new_n821), .B2(new_n667), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n825), .A2(new_n606), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(KEYINPUT109), .A3(new_n823), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n806), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n679), .A2(new_n743), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n840), .A2(new_n849), .ZN(new_n856));
  INV_X1    g670(.A(new_n806), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n806), .A2(new_n826), .A3(new_n839), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n857), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n862), .B2(new_n853), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n730), .A2(new_n751), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n776), .A2(new_n870), .A3(new_n371), .A4(new_n778), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n776), .A2(new_n371), .A3(new_n778), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT110), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n868), .A2(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n749), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT48), .Z(new_n876));
  AOI21_X1  g690(.A(new_n737), .B1(new_n873), .B2(new_n871), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n730), .A3(new_n702), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT118), .Z(new_n879));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n316), .A2(G952), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n745), .A2(new_n695), .A3(new_n370), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n868), .B2(new_n869), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n883), .B2(new_n704), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n880), .B1(new_n879), .B2(new_n884), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n876), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n797), .A2(new_n416), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n790), .B2(new_n792), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n891));
  INV_X1    g705(.A(new_n877), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n772), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT51), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n874), .A2(new_n742), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n367), .A2(new_n634), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n883), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n691), .A2(new_n313), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n877), .A2(new_n730), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT112), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT50), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n877), .A2(KEYINPUT112), .A3(new_n730), .A4(new_n901), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT50), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n900), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n896), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n912), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  INV_X1    g730(.A(new_n895), .ZN(new_n917));
  INV_X1    g731(.A(new_n893), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n890), .B2(KEYINPUT116), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT117), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n887), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n790), .A2(new_n792), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(KEYINPUT111), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n889), .B1(new_n923), .B2(KEYINPUT111), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n916), .B1(new_n912), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT115), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT115), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n916), .C1(new_n912), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n866), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(G952), .A2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n802), .B1(new_n932), .B2(new_n933), .ZN(G75));
  NOR3_X1   g748(.A1(new_n826), .A2(new_n860), .A3(new_n839), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n857), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n850), .B2(KEYINPUT53), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(G210), .A3(G902), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n303), .A2(new_n304), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n212), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n305), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n316), .A2(G952), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT121), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT120), .B1(new_n863), .B2(new_n285), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n937), .A2(new_n950), .A3(G902), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n188), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n944), .A2(KEYINPUT56), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(G51));
  XNOR2_X1  g768(.A(new_n937), .B(new_n864), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n765), .B(KEYINPUT57), .Z(new_n956));
  OAI21_X1  g770(.A(new_n467), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n949), .A2(new_n764), .A3(new_n951), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n946), .B1(new_n957), .B2(new_n958), .ZN(G54));
  AND2_X1   g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n949), .A2(new_n951), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n361), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n946), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n949), .A2(new_n361), .A3(new_n951), .A4(new_n960), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G60));
  AND2_X1   g780(.A1(new_n627), .A2(new_n629), .ZN(new_n967));
  XNOR2_X1  g781(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n410), .A2(new_n285), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n947), .B1(new_n955), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n967), .B1(new_n866), .B2(new_n970), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT60), .Z(new_n976));
  OAI211_X1 g790(.A(new_n659), .B(new_n976), .C1(new_n858), .C2(new_n861), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n937), .A2(new_n979), .A3(new_n659), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n601), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n937), .B2(new_n976), .ZN(new_n983));
  INV_X1    g797(.A(new_n947), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n985), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n984), .B(new_n983), .C1(new_n978), .C2(new_n980), .ZN(new_n987));
  XOR2_X1   g801(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(G66));
  INV_X1    g803(.A(new_n372), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n316), .B1(new_n990), .B2(G224), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n826), .A2(new_n844), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n316), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n941), .B1(G898), .B2(new_n316), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(G69));
  AND2_X1   g809(.A1(new_n351), .A2(new_n352), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n520), .B(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(G900), .B2(G953), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n783), .A2(new_n794), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n679), .A2(new_n712), .A3(new_n743), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n733), .A2(new_n749), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n832), .B1(new_n771), .B2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n999), .B1(new_n1004), .B2(new_n316), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1000), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1001), .A2(new_n700), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n635), .B1(new_n412), .B2(new_n367), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT125), .ZN(new_n1013));
  OR4_X1    g827(.A1(new_n604), .A2(new_n684), .A3(new_n750), .A4(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1015), .A2(new_n316), .ZN(new_n1016));
  INV_X1    g830(.A(new_n997), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1006), .B(new_n1007), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1015), .B2(new_n316), .ZN(new_n1019));
  OAI21_X1  g833(.A(KEYINPUT126), .B1(new_n1019), .B2(new_n1005), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n316), .B1(G227), .B2(G900), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1021), .ZN(new_n1023));
  OAI211_X1 g837(.A(KEYINPUT126), .B(new_n1023), .C1(new_n1019), .C2(new_n1005), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1022), .A2(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n1004), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n992), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n521), .A3(new_n553), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1027), .B1(new_n1015), .B2(new_n992), .ZN(new_n1031));
  INV_X1    g845(.A(new_n553), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1031), .A2(new_n486), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1030), .A2(new_n1033), .A3(new_n964), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n855), .A2(new_n858), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1027), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1032), .A2(new_n521), .ZN(new_n1037));
  OR2_X1    g851(.A1(new_n1037), .A2(KEYINPUT127), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n692), .B1(new_n1037), .B2(KEYINPUT127), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1034), .B1(new_n1035), .B2(new_n1040), .ZN(G57));
endmodule


