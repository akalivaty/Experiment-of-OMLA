//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n203), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n219), .A2(new_n220), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n214), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT68), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n214), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT66), .B(KEYINPUT0), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G20), .ZN(new_n235));
  OAI21_X1  g0035(.A(G50), .B1(G58), .B2(G68), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n232), .B1(new_n235), .B2(new_n236), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n228), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT70), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  AOI21_X1  g0056(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(G1), .B(G13), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n259), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(G226), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT71), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n261), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(KEYINPUT71), .A3(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G222), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G223), .A3(G1698), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n277), .B(new_n278), .C1(new_n203), .C2(new_n275), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n260), .B(new_n266), .C1(new_n279), .C2(new_n257), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n234), .B1(new_n213), .B2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n202), .A2(new_n212), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n212), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n284), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n211), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(new_n296), .B2(new_n294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n280), .B2(G169), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n282), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n299), .B(KEYINPUT9), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n280), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n280), .A2(G190), .ZN(new_n305));
  OR3_X1    g0105(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT10), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n275), .A2(G226), .A3(new_n276), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n275), .A2(G232), .A3(G1698), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G97), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n257), .ZN(new_n313));
  INV_X1    g0113(.A(new_n260), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(new_n217), .B2(new_n264), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(G190), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n313), .B2(new_n316), .ZN(new_n322));
  AOI211_X1 g0122(.A(KEYINPUT13), .B(new_n315), .C1(new_n312), .C2(new_n257), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n211), .A2(G20), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n295), .A2(G68), .A3(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n203), .B2(new_n287), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n284), .A2(new_n328), .A3(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n294), .A2(new_n216), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT11), .B1(new_n284), .B2(new_n328), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n321), .A2(new_n324), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n322), .A2(new_n323), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT14), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n318), .A2(G179), .A3(new_n320), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(G169), .C1(new_n322), .C2(new_n323), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n334), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(G223), .A2(G1698), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G226), .B2(new_n276), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n268), .A2(new_n269), .ZN(new_n348));
  INV_X1    g0148(.A(G87), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n347), .A2(new_n348), .B1(new_n261), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n257), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n260), .B1(G232), .B2(new_n265), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(KEYINPUT75), .A3(new_n257), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n353), .A2(new_n281), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n351), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n338), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G58), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n216), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(G20), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(G159), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n364), .B(new_n366), .C1(new_n367), .C2(new_n290), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n272), .A2(new_n273), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G20), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n348), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n216), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT16), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n270), .B2(new_n274), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n368), .B1(G68), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n375), .B(new_n284), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n286), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n325), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n295), .A2(new_n383), .B1(new_n294), .B2(new_n286), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n359), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n387));
  INV_X1    g0187(.A(G190), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n353), .A2(new_n388), .A3(new_n354), .A4(new_n355), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n357), .A2(new_n303), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n380), .A2(new_n391), .A3(new_n384), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n387), .A2(new_n394), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n286), .A2(new_n290), .B1(new_n212), .B2(new_n203), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n287), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n284), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n203), .B1(new_n211), .B2(G20), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n295), .A2(new_n407), .B1(new_n203), .B2(new_n294), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n314), .B1(new_n218), .B2(new_n264), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(new_n206), .C2(new_n275), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(new_n257), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G190), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n410), .B(new_n416), .C1(new_n303), .C2(new_n415), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n281), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n409), .C1(G169), .C2(new_n415), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n308), .A2(new_n345), .A3(new_n400), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G250), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n276), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n270), .A2(new_n274), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT76), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n270), .A2(new_n274), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(G244), .B(new_n276), .C1(new_n268), .C2(new_n269), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n270), .A2(new_n274), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n431), .B(new_n432), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n257), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT77), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n257), .C1(new_n428), .C2(new_n435), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(G257), .A3(new_n263), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(new_n263), .A3(G274), .A4(new_n441), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n445), .B2(new_n447), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n450), .A2(new_n451), .A3(G179), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n437), .A2(new_n439), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n293), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n211), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n283), .A2(new_n293), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(G97), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT6), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n459), .A2(new_n205), .A3(G107), .ZN(new_n460));
  XNOR2_X1  g0260(.A(G97), .B(G107), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n462), .A2(new_n212), .B1(new_n203), .B2(new_n290), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n377), .B2(G107), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n458), .B1(new_n464), .B2(new_n283), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n450), .A2(new_n451), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n436), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n338), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n453), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT79), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n377), .A2(G107), .ZN(new_n472));
  INV_X1    g0272(.A(new_n463), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n284), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n475), .A2(new_n458), .B1(new_n467), .B2(new_n338), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT79), .B1(new_n476), .B2(new_n453), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NOR4_X1   g0278(.A1(new_n257), .A2(KEYINPUT80), .A3(new_n441), .A4(new_n422), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n441), .A2(new_n422), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n263), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n263), .A2(G274), .A3(new_n441), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G116), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G238), .A2(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n218), .B2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n370), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n484), .B1(new_n489), .B2(new_n263), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n281), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT19), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n212), .B1(new_n311), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G87), .B2(new_n207), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n287), .B2(new_n205), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n370), .A2(new_n212), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n216), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(new_n284), .B1(new_n294), .B2(new_n402), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n402), .B2(new_n456), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n338), .B1(new_n483), .B2(new_n490), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n492), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n483), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n489), .A2(new_n263), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(G190), .A3(new_n504), .A4(new_n484), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n457), .A2(KEYINPUT81), .A3(G87), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT81), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n456), .B2(new_n349), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G200), .B1(new_n483), .B2(new_n490), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n499), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n437), .A2(new_n439), .A3(new_n466), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n436), .A2(new_n466), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n465), .B1(new_n515), .B2(G190), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n478), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT86), .ZN(new_n519));
  AOI21_X1  g0319(.A(G1698), .B1(new_n272), .B2(new_n273), .ZN(new_n520));
  AND2_X1   g0320(.A1(G257), .A2(G1698), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n268), .B2(new_n269), .ZN(new_n522));
  AOI22_X1  g0322(.A1(G250), .A2(new_n520), .B1(new_n522), .B2(KEYINPUT84), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n261), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G257), .A2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n272), .B2(new_n273), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT85), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(new_n276), .C1(new_n268), .C2(new_n269), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n527), .B2(new_n528), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n528), .B(new_n521), .C1(new_n268), .C2(new_n269), .ZN(new_n533));
  INV_X1    g0333(.A(new_n525), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n519), .B(new_n257), .C1(new_n530), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n257), .B1(new_n441), .B2(new_n446), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G264), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n447), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n536), .B1(new_n532), .B2(new_n535), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n529), .A2(KEYINPUT85), .A3(new_n545), .A4(new_n531), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n519), .B1(new_n547), .B2(new_n257), .ZN(new_n548));
  OAI21_X1  g0348(.A(G169), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n263), .B1(new_n544), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n541), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G179), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT25), .ZN(new_n555));
  AOI211_X1 g0355(.A(G107), .B(new_n293), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n457), .B2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT22), .B1(new_n497), .B2(new_n349), .ZN(new_n562));
  OR3_X1    g0362(.A1(new_n349), .A2(KEYINPUT22), .A3(G20), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n433), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n212), .A2(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n565), .B(KEYINPUT23), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n485), .B2(G20), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n486), .A2(KEYINPUT82), .A3(new_n212), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n564), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n561), .B1(new_n575), .B2(new_n284), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n553), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n543), .A2(G190), .A3(new_n548), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n551), .A2(G200), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n457), .A2(G116), .ZN(new_n583));
  INV_X1    g0383(.A(G116), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n294), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n212), .A2(G116), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n283), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n432), .B(new_n212), .C1(G33), .C2(new_n205), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n587), .A2(KEYINPUT20), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT20), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n583), .B(new_n585), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n276), .A2(G264), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n370), .B(new_n592), .C1(G257), .C2(G1698), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n275), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n257), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n539), .A2(G270), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(new_n447), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n591), .A2(new_n599), .A3(G169), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n599), .A2(new_n281), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n591), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n591), .A2(new_n599), .A3(KEYINPUT21), .A4(G169), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n599), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n591), .B1(G200), .B2(new_n599), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n582), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n421), .A2(new_n518), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT87), .ZN(G372));
  INV_X1    g0413(.A(new_n421), .ZN(new_n614));
  INV_X1    g0414(.A(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n578), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(new_n478), .A3(new_n517), .A4(new_n581), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT26), .B1(new_n478), .B2(new_n512), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n469), .A2(new_n512), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n617), .A2(new_n618), .A3(new_n502), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT88), .Z(new_n624));
  XNOR2_X1  g0424(.A(new_n392), .B(KEYINPUT17), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n335), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n318), .A2(new_n320), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n341), .B1(new_n627), .B2(G169), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n342), .A2(new_n340), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n344), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n626), .B1(new_n630), .B2(new_n419), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n385), .B(KEYINPUT18), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n307), .B2(new_n306), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n301), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n624), .A2(new_n636), .ZN(G369));
  NAND3_X1  g0437(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT89), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n591), .ZN(new_n645));
  MUX2_X1   g0445(.A(new_n610), .B(new_n606), .S(new_n645), .Z(new_n646));
  XNOR2_X1  g0446(.A(KEYINPUT90), .B(G330), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT91), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n644), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n582), .B1(new_n576), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n578), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n644), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n615), .A2(new_n644), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n582), .A2(new_n659), .B1(new_n654), .B2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n229), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT92), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n666), .A2(new_n667), .B1(new_n236), .B2(new_n664), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n667), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT93), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT28), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n622), .A2(new_n652), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT29), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n469), .A2(new_n470), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n476), .A2(KEYINPUT79), .A3(new_n453), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n512), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n620), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n620), .B2(new_n619), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n517), .A2(new_n581), .A3(new_n674), .A4(new_n675), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n606), .B1(new_n553), .B2(new_n577), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n502), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n652), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n491), .A2(new_n540), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n686), .A2(new_n599), .A3(new_n281), .ZN(new_n687));
  INV_X1    g0487(.A(new_n550), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n515), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n607), .A2(new_n491), .A3(G179), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n692), .B(new_n513), .C1(new_n550), .C2(new_n541), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n687), .A2(KEYINPUT30), .A3(new_n515), .A4(new_n688), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n644), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n611), .A2(new_n518), .A3(new_n644), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n648), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n685), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n671), .B1(new_n704), .B2(G1), .ZN(G364));
  INV_X1    g0505(.A(G13), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G45), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n663), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n233), .B1(G20), .B2(new_n338), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n212), .A2(new_n281), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n388), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G326), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n717), .A2(G190), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OR2_X1    g0523(.A1(KEYINPUT33), .A2(G317), .ZN(new_n724));
  NAND2_X1  g0524(.A1(KEYINPUT33), .A2(G317), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n281), .A2(new_n303), .A3(G190), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n721), .B(new_n726), .C1(G294), .C2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n212), .A2(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G190), .A3(G200), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G303), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G190), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n716), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n730), .A2(new_n737), .ZN(new_n740));
  INV_X1    g0540(.A(G329), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n716), .A2(G190), .A3(new_n303), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(G322), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n730), .A2(new_n388), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n275), .B1(G283), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n729), .A2(new_n736), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n206), .ZN(new_n750));
  INV_X1    g0550(.A(new_n728), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n723), .A2(new_n216), .B1(new_n205), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n750), .B(new_n752), .C1(G50), .C2(new_n718), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n735), .A2(G87), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT96), .B(G159), .Z(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n740), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n743), .A2(new_n360), .B1(new_n738), .B2(new_n203), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n433), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n753), .A2(new_n754), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n715), .B1(new_n749), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n714), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n662), .A2(new_n370), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n236), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n255), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n275), .A2(new_n229), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n209), .A2(new_n769), .B1(G116), .B2(new_n229), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n713), .B(new_n761), .C1(new_n765), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n764), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n646), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n713), .B1(new_n646), .B2(new_n648), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n651), .B2(new_n775), .ZN(G396));
  OAI21_X1  g0576(.A(KEYINPUT98), .B1(new_n419), .B2(new_n652), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n415), .A2(G169), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n410), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT98), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n779), .A2(new_n780), .A3(new_n418), .A4(new_n644), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n419), .B(new_n417), .C1(new_n410), .C2(new_n652), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT99), .Z(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(new_n672), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n644), .B1(new_n782), .B2(new_n783), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n621), .B1(new_n676), .B2(new_n620), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n681), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT101), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(KEYINPUT101), .B(new_n787), .C1(new_n681), .C2(new_n788), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n786), .A2(KEYINPUT100), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(KEYINPUT100), .B2(new_n786), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n702), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT102), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n712), .B1(new_n794), .B2(new_n702), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n714), .A2(new_n762), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n713), .B1(new_n203), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n755), .ZN(new_n801));
  INV_X1    g0601(.A(new_n738), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n744), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n719), .C1(new_n288), .C2(new_n723), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n734), .A2(new_n296), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n751), .A2(new_n360), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n370), .B1(new_n740), .B2(new_n810), .C1(new_n216), .C2(new_n746), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n805), .A2(new_n806), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n735), .A2(G107), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n815), .A2(new_n723), .B1(new_n719), .B2(new_n594), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G87), .B2(new_n747), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n743), .A2(new_n524), .B1(new_n740), .B2(new_n739), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G116), .B2(new_n802), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n275), .B1(G97), .B2(new_n728), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n784), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n800), .B1(new_n822), .B2(new_n715), .C1(new_n823), .C2(new_n763), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n798), .A2(new_n824), .ZN(G384));
  INV_X1    g0625(.A(new_n462), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n584), .B(new_n235), .C1(new_n826), .C2(KEYINPUT35), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(KEYINPUT35), .B2(new_n826), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  OAI21_X1  g0629(.A(G77), .B1(new_n360), .B2(new_n216), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(new_n236), .B1(G50), .B2(new_n216), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(G1), .A3(new_n706), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT103), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n684), .A2(new_n614), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n636), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT108), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT109), .ZN(new_n838));
  INV_X1    g0638(.A(new_n384), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n284), .B1(new_n374), .B2(new_n379), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(KEYINPUT105), .B1(KEYINPUT16), .B2(new_n374), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT105), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n284), .C1(new_n374), .C2(new_n379), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n392), .B1(new_n844), .B2(new_n359), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n642), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT37), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n393), .A2(new_n385), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n380), .A2(new_n384), .ZN(new_n849));
  INV_X1    g0649(.A(new_n642), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT37), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n399), .A2(new_n846), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n344), .A2(new_n644), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n630), .A2(new_n335), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n344), .B(new_n644), .C1(new_n343), .C2(new_n336), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n791), .A2(new_n792), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n419), .A2(new_n644), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(KEYINPUT104), .B(new_n865), .C1(new_n791), .C2(new_n792), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n858), .B(new_n862), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n633), .A2(new_n642), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT106), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n849), .A2(new_n850), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n386), .A2(new_n875), .A3(new_n392), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n848), .A2(new_n876), .A3(KEYINPUT37), .A4(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n875), .B1(new_n632), .B2(new_n625), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n874), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT39), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(KEYINPUT39), .B2(new_n857), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n343), .A2(new_n344), .A3(new_n652), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n869), .A2(KEYINPUT106), .A3(new_n870), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n873), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n838), .B(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n478), .A2(new_n517), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n610), .A3(new_n582), .A4(new_n652), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n895), .A2(KEYINPUT111), .B1(new_n696), .B2(new_n699), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT111), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n695), .A2(new_n897), .A3(KEYINPUT31), .A4(new_n644), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n784), .B1(new_n860), .B2(new_n861), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n899), .B(new_n900), .C1(new_n855), .C2(new_n856), .ZN(new_n901));
  XNOR2_X1  g0701(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n862), .A2(new_n823), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n895), .A2(KEYINPUT111), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n696), .A2(new_n699), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n903), .B1(new_n907), .B2(new_n894), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n883), .B2(new_n884), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n901), .A2(new_n902), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n899), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n421), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n614), .A3(new_n899), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n648), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n892), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n211), .B2(new_n707), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n892), .A2(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n834), .B1(new_n918), .B2(new_n919), .ZN(G367));
  AOI22_X1  g0720(.A1(new_n514), .A2(new_n516), .B1(new_n465), .B2(new_n644), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n478), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n476), .A2(new_n453), .A3(new_n644), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n582), .A2(new_n659), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT112), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n477), .B(new_n471), .C1(new_n924), .C2(new_n654), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n930), .C1(new_n644), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n509), .A2(new_n499), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n644), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n502), .A3(new_n511), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n502), .B2(new_n934), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n932), .A2(KEYINPUT43), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n932), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n658), .B2(new_n925), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n658), .A2(new_n925), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n663), .B(KEYINPUT41), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n926), .B1(new_n657), .B2(new_n659), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n650), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n703), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n660), .A2(new_n924), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT45), .Z(new_n953));
  NOR2_X1   g0753(.A1(new_n660), .A2(new_n924), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n658), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n951), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n946), .B1(new_n958), .B2(new_n704), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n943), .B(new_n945), .C1(new_n711), .C2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n766), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n765), .B1(new_n229), .B2(new_n402), .C1(new_n961), .C2(new_n248), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(new_n712), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n723), .A2(new_n755), .B1(new_n216), .B2(new_n751), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G143), .B2(new_n718), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n735), .A2(G58), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n738), .A2(new_n296), .B1(new_n740), .B2(new_n804), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G150), .B2(new_n744), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n433), .B1(G77), .B2(new_n747), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n965), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n718), .A2(G311), .B1(G107), .B2(new_n728), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n743), .A2(new_n594), .B1(new_n738), .B2(new_n815), .ZN(new_n972));
  INV_X1    g0772(.A(new_n740), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n370), .B(new_n972), .C1(G317), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n735), .A2(KEYINPUT46), .A3(G116), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n722), .A2(G294), .B1(new_n747), .B2(G97), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT46), .B1(new_n735), .B2(G116), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n970), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  OAI221_X1 g0780(.A(new_n963), .B1(new_n773), .B2(new_n936), .C1(new_n980), .C2(new_n715), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n960), .A2(new_n981), .ZN(G387));
  NAND2_X1  g0782(.A1(new_n950), .A2(new_n951), .ZN(new_n983));
  INV_X1    g0783(.A(new_n948), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n663), .C1(new_n704), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n656), .A2(new_n764), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n243), .A2(G45), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n987), .A2(new_n961), .B1(new_n665), .B2(new_n769), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n286), .B2(G50), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n381), .A2(new_n989), .A3(new_n296), .ZN(new_n992));
  AOI21_X1  g0792(.A(G45), .B1(G68), .B2(G77), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(new_n665), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n988), .A2(new_n994), .B1(new_n206), .B2(new_n662), .ZN(new_n995));
  INV_X1    g0795(.A(new_n765), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n712), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n743), .A2(new_n296), .B1(new_n740), .B2(new_n288), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n348), .B(new_n998), .C1(G68), .C2(new_n802), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n735), .A2(G77), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n751), .A2(new_n402), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G97), .B2(new_n747), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G159), .A2(new_n718), .B1(new_n722), .B2(new_n381), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n370), .B1(new_n973), .B2(G326), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n743), .A2(new_n1006), .B1(new_n738), .B2(new_n594), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT115), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(KEYINPUT115), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G311), .A2(new_n722), .B1(new_n718), .B2(G322), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n735), .A2(G294), .B1(G283), .B2(new_n728), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT49), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT116), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1005), .B1(new_n584), .B2(new_n746), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1017), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(KEYINPUT116), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1004), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n997), .B1(new_n1022), .B2(new_n714), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n984), .A2(new_n711), .B1(new_n986), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n985), .A2(new_n1024), .ZN(G393));
  INV_X1    g0825(.A(new_n957), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n983), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1027), .A2(new_n663), .A3(new_n958), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n766), .A2(new_n252), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n765), .C1(new_n205), .C2(new_n229), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n751), .A2(new_n203), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n381), .B2(new_n802), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n296), .B2(new_n723), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT118), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G150), .A2(new_n718), .B1(new_n744), .B2(G159), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n370), .B1(new_n746), .B2(new_n349), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n735), .A2(G68), .B1(G143), .B2(new_n973), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT117), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n719), .A2(new_n1006), .B1(new_n739), .B2(new_n743), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n751), .A2(new_n584), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n750), .B(new_n1045), .C1(G303), .C2(new_n722), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n738), .A2(new_n524), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G322), .B2(new_n973), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n433), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G283), .B2(new_n735), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1040), .A2(new_n1042), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n712), .B(new_n1030), .C1(new_n1051), .C2(new_n715), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n925), .B2(new_n764), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n957), .B2(new_n711), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1028), .A2(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n883), .A2(new_n884), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n682), .A2(new_n784), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1057), .A2(new_n866), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n862), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n887), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT101), .B1(new_n622), .B2(new_n787), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n792), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n866), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT104), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n864), .A2(new_n863), .A3(new_n866), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n888), .B1(new_n1066), .B2(new_n862), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1060), .B1(new_n1067), .B2(new_n886), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n899), .A2(G330), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n900), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n702), .A2(new_n784), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n862), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1060), .B(new_n1075), .C1(new_n1067), .C2(new_n886), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n835), .B(new_n636), .C1(new_n421), .C2(new_n1069), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1071), .B1(new_n1074), .B2(new_n862), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1066), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1059), .B1(new_n1069), .B2(new_n785), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1075), .A2(new_n1058), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1078), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1073), .A2(new_n1076), .A3(new_n1083), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n663), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1073), .A2(new_n1076), .A3(new_n711), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n713), .B1(new_n286), .B2(new_n799), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n719), .A2(new_n815), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1031), .B(new_n1090), .C1(G107), .C2(new_n722), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n738), .A2(new_n205), .B1(new_n740), .B2(new_n524), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G116), .B2(new_n744), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n275), .B1(G68), .B2(new_n747), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n754), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n744), .A2(G132), .B1(new_n973), .B2(G125), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT54), .B(G143), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n738), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n433), .B(new_n1098), .C1(G128), .C2(new_n718), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT53), .B1(new_n734), .B2(new_n288), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n723), .A2(new_n804), .B1(new_n367), .B2(new_n751), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G50), .B2(new_n747), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n734), .A2(KEYINPUT53), .A3(new_n288), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1095), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT119), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n714), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1089), .B1(new_n1107), .B2(new_n1109), .C1(new_n886), .C2(new_n763), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1087), .A2(new_n1111), .ZN(G378));
  XNOR2_X1  g0912(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n850), .A2(new_n299), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n308), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n308), .A2(new_n1115), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1118), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n1116), .A3(new_n1113), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n911), .B2(G330), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n900), .B1(new_n906), .B2(new_n701), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n902), .B1(new_n857), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n908), .A2(new_n910), .ZN(new_n1126));
  AND4_X1   g0926(.A1(G330), .A2(new_n1125), .A3(new_n1126), .A4(new_n1122), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n890), .A2(new_n889), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT106), .B1(new_n869), .B2(new_n870), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n891), .A2(KEYINPUT121), .A3(new_n1129), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT122), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n1128), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n873), .A2(new_n889), .A3(new_n1128), .A4(new_n890), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(KEYINPUT122), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1134), .B(new_n1135), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1078), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1086), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT57), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(KEYINPUT57), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n663), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n744), .A2(G128), .B1(new_n802), .B2(G137), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n810), .B2(new_n723), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n718), .A2(G125), .B1(G150), .B2(new_n728), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT120), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1097), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1150), .B(new_n1152), .C1(new_n735), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT59), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n801), .A2(new_n747), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n973), .C2(G124), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n296), .B1(G33), .B2(G41), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n348), .B2(new_n262), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n743), .A2(new_n206), .B1(new_n738), .B2(new_n402), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n348), .B(new_n262), .C1(new_n740), .C2(new_n815), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n746), .A2(new_n360), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G68), .B2(new_n728), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G97), .A2(new_n722), .B1(new_n718), .B2(G116), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1000), .A2(new_n1165), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT58), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1162), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1160), .B(new_n1171), .C1(new_n1170), .C2(new_n1169), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n714), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n713), .B1(new_n296), .B2(new_n799), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n1122), .C2(new_n763), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1141), .B2(new_n711), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1148), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G375));
  NAND2_X1  g0980(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1078), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n946), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1084), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n723), .A2(new_n584), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1001), .B(new_n1186), .C1(G294), .C2(new_n718), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n735), .A2(G97), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n738), .A2(new_n206), .B1(new_n740), .B2(new_n594), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G283), .B2(new_n744), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n275), .B1(G77), .B2(new_n747), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n743), .A2(new_n804), .B1(new_n738), .B2(new_n288), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n348), .B(new_n1193), .C1(G128), .C2(new_n973), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n735), .A2(G159), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1166), .B1(G50), .B2(new_n728), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G132), .A2(new_n718), .B1(new_n722), .B2(new_n1153), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n715), .B1(new_n1192), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n713), .B(new_n1199), .C1(new_n216), .C2(new_n799), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT123), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n763), .B2(new_n862), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n711), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1182), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1185), .A2(new_n1205), .ZN(G381));
  OR3_X1    g1006(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1207), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1208));
  INV_X1    g1008(.A(G378), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n1179), .ZN(G407));
  NAND4_X1  g1010(.A1(new_n1179), .A2(G213), .A3(new_n643), .A4(new_n1209), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(G407), .A2(G213), .A3(new_n1211), .ZN(G409));
  OAI211_X1 g1012(.A(G378), .B(new_n1177), .C1(new_n1144), .C2(new_n1147), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1139), .B(new_n1136), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1184), .B(new_n1143), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1176), .B1(new_n1145), .B2(new_n711), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1209), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1213), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT124), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n643), .A2(G213), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1213), .A2(new_n1219), .A3(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n798), .A2(new_n824), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1183), .B1(new_n1226), .B2(new_n1083), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1182), .A2(KEYINPUT60), .A3(new_n1078), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n663), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1205), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1225), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G384), .A2(new_n1205), .A3(new_n1229), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT63), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n960), .A2(new_n981), .A3(G390), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(G396), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G390), .B1(new_n960), .B2(new_n981), .ZN(new_n1241));
  OR3_X1    g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT61), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n643), .A2(G213), .A3(G2897), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1231), .A2(new_n1232), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1247), .A2(new_n1248), .A3(KEYINPUT125), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1224), .A2(new_n1222), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1223), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1251), .A2(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1234), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1237), .A2(new_n1245), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1256), .B2(new_n1249), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1235), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1256), .A2(KEYINPUT62), .A3(new_n1234), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1260), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1244), .B(KEYINPUT126), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1258), .B1(new_n1264), .B2(new_n1265), .ZN(G405));
  NAND2_X1  g1066(.A1(G375), .A2(new_n1209), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1213), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1234), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1213), .A3(new_n1233), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1244), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1242), .A3(new_n1243), .A4(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(G402));
endmodule


