//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g0008(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n218), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n221), .B1(KEYINPUT1), .B2(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n214), .B(new_n229), .C1(KEYINPUT1), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G223), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n252), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G222), .A3(new_n248), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n254), .B(new_n256), .C1(new_n257), .C2(new_n255), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n210), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(new_n215), .C1(G41), .C2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n206), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n268), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n265), .B1(new_n270), .B2(G226), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G169), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G58), .ZN(new_n279));
  INV_X1    g0079(.A(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT8), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT69), .ZN(new_n282));
  OR3_X1    g0082(.A1(new_n280), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n216), .A2(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n208), .A2(new_n209), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n288), .B1(new_n202), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n215), .A2(G20), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n208), .A2(new_n289), .A3(new_n209), .A4(new_n287), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n294), .ZN(new_n296));
  OAI211_X1 g0096(.A(G50), .B(new_n292), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n275), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n291), .B2(new_n297), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n272), .A2(G190), .ZN(new_n303));
  AOI21_X1  g0103(.A(G200), .B1(new_n262), .B2(new_n271), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n300), .A2(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n298), .B(KEYINPUT9), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n272), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G190), .B2(new_n272), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n306), .A3(KEYINPUT10), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT71), .ZN(new_n316));
  INV_X1    g0116(.A(new_n276), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n319), .A2(new_n285), .B1(new_n216), .B2(new_n257), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n288), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n293), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n292), .ZN(new_n323));
  MUX2_X1   g0123(.A(new_n289), .B(new_n323), .S(G77), .Z(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n253), .A2(G238), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n255), .A2(G232), .A3(new_n248), .ZN(new_n327));
  INV_X1    g0127(.A(G107), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n255), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n261), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n265), .B1(new_n270), .B2(G244), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n332), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n311), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n325), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(G169), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(G179), .A3(new_n332), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n338), .B1(new_n321), .B2(new_n324), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  AND4_X1   g0140(.A1(new_n299), .A2(new_n309), .A3(new_n314), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n215), .A2(G13), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G68), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(G20), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n344), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n257), .B2(new_n285), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n288), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n350), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n344), .B2(new_n323), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n265), .B1(new_n270), .B2(G238), .ZN(new_n354));
  AND2_X1   g0154(.A1(KEYINPUT3), .A2(G33), .ZN(new_n355));
  NOR2_X1   g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  OAI211_X1 g0156(.A(G232), .B(G1698), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(G226), .B(new_n248), .C1(new_n355), .C2(new_n356), .ZN(new_n358));
  AND3_X1   g0158(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT74), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n261), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n261), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n354), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT13), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n354), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(G179), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n369), .ZN(new_n372));
  AND2_X1   g0172(.A1(KEYINPUT75), .A2(G169), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n370), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n372), .A2(new_n371), .A3(new_n373), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n353), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n311), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n367), .A2(new_n331), .A3(new_n369), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n353), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n341), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n282), .A2(new_n283), .A3(new_n292), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n295), .B2(new_n296), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n284), .A2(new_n290), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n251), .A2(new_n216), .A3(new_n252), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n252), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n344), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n280), .A2(new_n344), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n393), .B2(new_n201), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n276), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT16), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n355), .A2(new_n356), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n398), .B2(new_n216), .ZN(new_n399));
  INV_X1    g0199(.A(new_n391), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n384), .A2(new_n386), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(new_n288), .B1(new_n406), .B2(KEYINPUT76), .ZN(new_n407));
  OAI211_X1 g0207(.A(G223), .B(new_n248), .C1(new_n355), .C2(new_n356), .ZN(new_n408));
  OAI211_X1 g0208(.A(G226), .B(G1698), .C1(new_n355), .C2(new_n356), .ZN(new_n409));
  INV_X1    g0209(.A(G87), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n250), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT77), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT77), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n408), .A2(new_n409), .A3(new_n415), .A4(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n261), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n265), .B1(new_n270), .B2(G232), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n331), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n266), .A2(new_n268), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n269), .A2(new_n259), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G232), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n265), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n416), .A2(new_n261), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n414), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n419), .B1(new_n426), .B2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n429));
  AND4_X1   g0229(.A1(new_n387), .A2(new_n407), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n208), .A2(new_n209), .A3(new_n287), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n397), .B2(new_n404), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n293), .A2(new_n294), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n382), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n386), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n434), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n432), .B1(new_n441), .B2(new_n427), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n430), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n402), .B1(new_n401), .B2(new_n403), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n392), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n288), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n406), .A2(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n387), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n411), .B1(new_n253), .B2(G226), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n415), .B1(new_n449), .B2(new_n408), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n416), .A2(new_n261), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n274), .B(new_n418), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(G169), .B1(new_n417), .B2(new_n418), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n448), .A2(new_n455), .A3(KEYINPUT18), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT18), .B1(new_n448), .B2(new_n455), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT78), .B(KEYINPUT18), .C1(new_n448), .C2(new_n455), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n443), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n381), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n250), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  AOI21_X1  g0264(.A(G20), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n216), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n288), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n289), .A2(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n215), .A2(G33), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT81), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n293), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G257), .B(new_n248), .C1(new_n355), .C2(new_n356), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n255), .A2(KEYINPUT84), .A3(G257), .A4(new_n248), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n253), .A2(G264), .B1(new_n398), .B2(G303), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n261), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT85), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n215), .A2(G45), .ZN(new_n487));
  OR2_X1    g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NAND2_X1  g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G274), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n421), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  INV_X1    g0293(.A(G270), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n485), .A2(new_n486), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n260), .B1(new_n482), .B2(new_n483), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT85), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n311), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(G190), .B1(new_n497), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n477), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  INV_X1    g0304(.A(G169), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n470), .B2(new_n475), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n497), .A3(new_n499), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n506), .A2(new_n497), .A3(KEYINPUT21), .A4(new_n499), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n498), .A2(new_n495), .A3(new_n274), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n476), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n486), .B1(new_n485), .B2(new_n496), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n498), .A2(new_n495), .A3(KEYINPUT85), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n331), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n500), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n477), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n504), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n216), .B(G87), .C1(new_n355), .C2(new_n356), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT22), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT23), .B1(new_n216), .B2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n466), .B2(new_n285), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n216), .A2(KEYINPUT23), .A3(G107), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n522), .A2(KEYINPUT24), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n288), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n343), .A2(G20), .A3(new_n328), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G107), .B2(new_n474), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n255), .A2(G250), .A3(new_n248), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n255), .A2(G257), .A3(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G294), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n261), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n490), .B1(new_n269), .B2(new_n259), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G264), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n491), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n540), .A2(new_n261), .B1(new_n542), .B2(G264), .ZN(new_n546));
  AOI21_X1  g0346(.A(G200), .B1(new_n546), .B2(new_n491), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n533), .B(new_n536), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G244), .B(G1698), .C1(new_n355), .C2(new_n356), .ZN(new_n549));
  OAI211_X1 g0349(.A(G238), .B(new_n248), .C1(new_n355), .C2(new_n356), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n250), .C2(new_n466), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n487), .A2(G250), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n264), .B2(new_n487), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n551), .A2(new_n261), .B1(new_n421), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n331), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G200), .B2(new_n554), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n255), .A2(new_n216), .A3(G68), .ZN(new_n557));
  INV_X1    g0357(.A(G97), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n250), .A2(new_n558), .A3(G20), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(KEYINPUT19), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT19), .B1(new_n359), .B2(new_n360), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G87), .A2(G97), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n216), .B1(new_n328), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n288), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n319), .A2(new_n290), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n474), .A2(G87), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n551), .A2(new_n261), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n553), .A2(new_n421), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(G179), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n505), .B2(new_n554), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n473), .A2(new_n293), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n564), .B(new_n565), .C1(new_n319), .C2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n556), .A2(new_n567), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n548), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(new_n248), .C1(new_n355), .C2(new_n356), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n576), .A2(new_n577), .B1(G33), .B2(G283), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n253), .A2(KEYINPUT82), .A3(G250), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT82), .B1(new_n253), .B2(G250), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n261), .ZN(new_n583));
  INV_X1    g0383(.A(G257), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n491), .B1(new_n493), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(KEYINPUT83), .A3(G200), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT83), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n585), .B1(new_n582), .B2(new_n261), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(new_n311), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n290), .A2(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n572), .B2(G97), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n317), .A2(new_n257), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  AND2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n328), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(KEYINPUT80), .B(new_n596), .C1(new_n602), .C2(new_n216), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n216), .B1(new_n600), .B2(new_n601), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n595), .ZN(new_n606));
  OAI21_X1  g0406(.A(G107), .B1(new_n399), .B2(new_n400), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n594), .B1(new_n608), .B2(new_n288), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n583), .A2(G190), .A3(new_n586), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n592), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n544), .A2(G169), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n274), .B2(new_n544), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n532), .A2(new_n288), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT24), .B1(new_n522), .B2(new_n528), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n536), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n608), .A2(new_n288), .ZN(new_n618));
  INV_X1    g0418(.A(new_n594), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n590), .A2(new_n505), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n274), .B(new_n585), .C1(new_n582), .C2(new_n261), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n575), .A2(new_n611), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n520), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n462), .A2(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n457), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n456), .ZN(new_n628));
  INV_X1    g0428(.A(new_n376), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n339), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n380), .A2(new_n443), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n309), .A2(new_n314), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n632), .A2(new_n633), .B1(new_n298), .B2(new_n275), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n509), .A2(new_n617), .A3(new_n510), .A4(new_n512), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(new_n575), .A3(new_n611), .A4(new_n623), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n556), .A2(new_n567), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n571), .A2(new_n573), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n623), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n587), .A2(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n590), .A2(G179), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n609), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n574), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n641), .A2(new_n646), .A3(new_n639), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n637), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n462), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n634), .A2(new_n649), .ZN(G369));
  OR3_X1    g0450(.A1(new_n342), .A2(KEYINPUT27), .A3(G20), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n342), .B2(G20), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n477), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n518), .B1(new_n517), .B2(new_n477), .ZN(new_n656));
  AOI211_X1 g0456(.A(KEYINPUT86), .B(new_n476), .C1(new_n516), .C2(new_n500), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n513), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n513), .B2(new_n655), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n617), .ZN(new_n663));
  INV_X1    g0463(.A(new_n654), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n616), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n548), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n654), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n513), .A2(new_n664), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n671), .A2(new_n668), .A3(new_n666), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n219), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G1), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n562), .A2(new_n328), .A3(new_n466), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT88), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n678), .A2(new_n680), .B1(new_n213), .B2(new_n677), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n587), .A2(new_n544), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n554), .A2(G179), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n497), .A2(new_n499), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT89), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT89), .A4(new_n684), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n546), .A2(new_n554), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n511), .A3(new_n590), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n690), .A2(new_n511), .A3(KEYINPUT30), .A4(new_n590), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n664), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n623), .A2(new_n548), .A3(new_n574), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n609), .A2(new_n610), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n591), .B2(new_n588), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n701), .A2(new_n703), .A3(new_n663), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n658), .A2(new_n704), .A3(new_n513), .A4(new_n654), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT31), .B(new_n664), .C1(new_n689), .C2(new_n695), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n696), .A2(KEYINPUT90), .A3(new_n697), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n700), .A2(new_n705), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n654), .B1(new_n637), .B2(new_n647), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n647), .A2(KEYINPUT91), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT91), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n641), .A2(new_n646), .A3(new_n715), .A4(new_n639), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n636), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT29), .B(new_n654), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n709), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n682), .B1(new_n719), .B2(G1), .ZN(G364));
  INV_X1    g0520(.A(G13), .ZN(new_n721));
  INV_X1    g0521(.A(G45), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(G20), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT92), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT92), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n676), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT93), .Z(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n210), .B1(new_n216), .B2(G169), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n216), .A2(G190), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G179), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G159), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n216), .A2(new_n331), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n274), .A2(new_n311), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n311), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G50), .A2(new_n740), .B1(new_n743), .B2(G107), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(new_n741), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n410), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n216), .B1(new_n732), .B2(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n558), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n738), .A2(new_n731), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n255), .B1(new_n749), .B2(new_n344), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n736), .A2(new_n746), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n274), .A2(G200), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT96), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n731), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n731), .B2(new_n752), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n737), .A2(new_n752), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n257), .B1(new_n280), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n751), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n739), .B(KEYINPUT98), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n756), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(G326), .B1(G311), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  INV_X1    g0566(.A(G329), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n757), .A2(new_n766), .B1(new_n733), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G294), .ZN(new_n769));
  INV_X1    g0569(.A(G303), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n398), .B1(new_n747), .B2(new_n769), .C1(new_n770), .C2(new_n745), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n768), .B(new_n771), .C1(G283), .C2(new_n743), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n749), .B1(new_n774), .B2(KEYINPUT99), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(KEYINPUT99), .B2(new_n774), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n765), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n730), .B1(new_n761), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n216), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n730), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT94), .Z(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT95), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n675), .A2(new_n398), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G355), .B1(new_n466), .B2(new_n675), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n675), .A2(new_n255), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n213), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n246), .A2(new_n722), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n729), .B(new_n778), .C1(new_n783), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT100), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n660), .B2(new_n780), .ZN(new_n792));
  INV_X1    g0592(.A(new_n727), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n661), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n660), .A2(G330), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT101), .Z(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  INV_X1    g0598(.A(KEYINPUT104), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n337), .A2(new_n338), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n325), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n801), .B2(new_n654), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n339), .A2(KEYINPUT104), .A3(new_n664), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n654), .B1(new_n321), .B2(new_n324), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n336), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT103), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n339), .A2(KEYINPUT103), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n804), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n710), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n709), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n727), .B1(new_n813), .B2(new_n709), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(new_n779), .ZN(new_n817));
  INV_X1    g0617(.A(new_n730), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n779), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n728), .B1(G77), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n749), .A2(KEYINPUT102), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n749), .A2(KEYINPUT102), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G283), .B1(G116), .B2(new_n764), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n742), .A2(new_n410), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n739), .A2(new_n770), .B1(new_n745), .B2(new_n328), .ZN(new_n827));
  INV_X1    g0627(.A(new_n757), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n826), .B(new_n827), .C1(G294), .C2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n255), .B(new_n748), .C1(G311), .C2(new_n734), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n255), .B1(new_n745), .B2(new_n202), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n742), .A2(new_n344), .B1(new_n733), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n747), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n834), .C1(G58), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n749), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G137), .A2(new_n740), .B1(new_n837), .B2(G150), .ZN(new_n838));
  INV_X1    g0638(.A(G143), .ZN(new_n839));
  INV_X1    g0639(.A(G159), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n839), .B2(new_n757), .C1(new_n756), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n836), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n831), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n821), .B1(new_n846), .B2(new_n818), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n815), .A2(new_n816), .B1(new_n817), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  XOR2_X1   g0649(.A(new_n602), .B(KEYINPUT35), .Z(new_n850));
  NOR3_X1   g0650(.A1(new_n850), .A2(new_n212), .A3(new_n466), .ZN(new_n851));
  XNOR2_X1  g0651(.A(KEYINPUT105), .B(KEYINPUT36), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OR3_X1    g0653(.A1(new_n393), .A2(new_n213), .A3(new_n257), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n202), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n215), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n628), .A2(new_n653), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n648), .A2(new_n654), .A3(new_n812), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n808), .A2(new_n809), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n654), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n372), .A2(new_n371), .A3(new_n373), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n370), .A2(new_n371), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n372), .A2(new_n373), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n353), .B(new_n664), .C1(new_n867), .C2(new_n379), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n353), .A2(new_n664), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n376), .A2(new_n380), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n446), .A2(new_n384), .A3(new_n386), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n653), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n461), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT106), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n461), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n448), .A2(new_n455), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT107), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n441), .A2(new_n427), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n448), .A2(new_n653), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n874), .B1(new_n455), .B2(new_n653), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n884), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n880), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n887), .B2(new_n888), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n452), .B1(new_n426), .B2(G169), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n407), .B2(new_n387), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT78), .B1(new_n899), .B2(KEYINPUT18), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n457), .A2(new_n458), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n456), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n875), .B1(new_n902), .B2(new_n443), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n897), .B1(new_n903), .B2(new_n879), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT108), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT38), .A4(new_n878), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n880), .A2(new_n894), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n879), .B1(new_n461), .B2(new_n876), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n896), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n858), .B1(new_n873), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n906), .A4(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n629), .A2(new_n654), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n908), .A2(new_n907), .A3(new_n909), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n886), .B2(new_n899), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n889), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n628), .A2(new_n443), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n448), .A3(new_n653), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n916), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n913), .A2(new_n915), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n718), .A2(new_n712), .A3(new_n462), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(new_n634), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n925), .B(new_n927), .Z(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n705), .A2(new_n706), .A3(new_n698), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n811), .B1(new_n868), .B2(new_n870), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n906), .A2(new_n910), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT40), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n917), .B2(new_n922), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT109), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n936), .B(KEYINPUT109), .C1(new_n917), .C2(new_n922), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n929), .A2(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n462), .A2(new_n930), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(G330), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(G1), .B1(new_n721), .B2(G20), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n928), .A2(new_n945), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n857), .B1(new_n948), .B2(new_n949), .ZN(G367));
  NAND2_X1  g0750(.A1(new_n644), .A2(new_n664), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT110), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n611), .B(new_n623), .C1(new_n609), .C2(new_n654), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n672), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT42), .Z(new_n956));
  NOR2_X1   g0756(.A1(new_n567), .A2(new_n654), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n574), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n639), .B2(new_n957), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n617), .B1(new_n952), .B2(new_n953), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n654), .B1(new_n961), .B2(new_n644), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n956), .A2(new_n962), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n959), .B(KEYINPUT43), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n670), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n954), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n970), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n676), .B(KEYINPUT41), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n673), .A2(new_n954), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT44), .B1(new_n673), .B2(new_n954), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n673), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n969), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n670), .A3(new_n977), .A4(new_n978), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n669), .B(new_n671), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n661), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n719), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n973), .B1(new_n986), .B2(new_n719), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n971), .B(new_n972), .C1(new_n726), .C2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n786), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n238), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n219), .A2(new_n319), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n990), .A2(new_n782), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n729), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n763), .A2(G311), .B1(G294), .B2(new_n824), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n745), .A2(new_n466), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G107), .B2(new_n835), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n764), .A2(G283), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n742), .A2(new_n558), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n398), .B1(new_n757), .B2(new_n770), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G317), .C2(new_n734), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n997), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n745), .A2(new_n280), .B1(new_n742), .B2(new_n257), .ZN(new_n1003));
  INV_X1    g0803(.A(G150), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n255), .B1(new_n747), .B2(new_n344), .C1(new_n757), .C2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G137), .C2(new_n734), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n824), .A2(G159), .B1(G50), .B2(new_n764), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n839), .C2(new_n762), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT47), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1002), .A2(new_n1008), .A3(KEYINPUT47), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n818), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n993), .B1(new_n1009), .B2(new_n1011), .C1(new_n959), .C2(new_n780), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n988), .A2(new_n1012), .ZN(G387));
  NOR2_X1   g0813(.A1(new_n985), .A2(new_n677), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n719), .B2(new_n983), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n983), .A2(new_n726), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n784), .A2(new_n680), .B1(new_n328), .B2(new_n675), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n680), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n316), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(KEYINPUT50), .B2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n786), .B1(new_n234), .B2(new_n722), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n729), .B1(new_n1024), .B2(new_n783), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n824), .A2(G311), .B1(G317), .B2(new_n828), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n770), .B2(new_n756), .C1(new_n766), .C2(new_n762), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  INV_X1    g0830(.A(G283), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n745), .A2(new_n769), .B1(new_n747), .B2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n398), .B1(new_n742), .B2(new_n466), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G326), .B2(new_n734), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n284), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n764), .A2(G68), .B1(new_n1039), .B2(new_n837), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n745), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G159), .A2(new_n740), .B1(new_n1041), .B2(G77), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G50), .A2(new_n828), .B1(new_n734), .B2(G150), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n747), .A2(new_n319), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n999), .A2(new_n1044), .A3(new_n398), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1025), .B1(new_n669), .B2(new_n780), .C1(new_n1047), .C2(new_n730), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1015), .A2(new_n1016), .A3(new_n1048), .ZN(G393));
  INV_X1    g0849(.A(new_n782), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n558), .B2(new_n219), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n243), .A2(new_n989), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n728), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G283), .A2(new_n1041), .B1(new_n734), .B2(G322), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n398), .C1(new_n328), .C2(new_n742), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G317), .A2(new_n740), .B1(new_n828), .B2(G311), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  INV_X1    g0857(.A(new_n824), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1057), .B1(new_n769), .B2(new_n756), .C1(new_n770), .C2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1055), .B(new_n1059), .C1(G116), .C2(new_n835), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n316), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n824), .A2(G50), .B1(new_n1064), .B2(new_n764), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n739), .A2(new_n1004), .B1(new_n757), .B2(new_n840), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n745), .A2(new_n344), .B1(new_n733), .B2(new_n839), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n747), .A2(new_n257), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1068), .A2(new_n826), .A3(new_n1069), .A4(new_n398), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1065), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1062), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1053), .B1(new_n1072), .B2(new_n818), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n780), .B2(new_n954), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n980), .A2(new_n981), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n726), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n986), .A2(new_n676), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n984), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(G390));
  OAI21_X1  g0881(.A(new_n728), .B1(new_n1039), .B2(new_n820), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n824), .A2(G107), .B1(G97), .B2(new_n764), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G68), .A2(new_n743), .B1(new_n734), .B2(G294), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G283), .A2(new_n740), .B1(new_n828), .B2(G116), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n255), .B(new_n1069), .C1(G87), .C2(new_n1041), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n745), .A2(new_n1004), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT53), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(KEYINPUT54), .B(G143), .ZN(new_n1090));
  INV_X1    g0890(.A(G137), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1089), .B1(new_n756), .B2(new_n1090), .C1(new_n1058), .C2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G128), .A2(new_n740), .B1(new_n743), .B2(G50), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n398), .B1(new_n734), .B2(G125), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n828), .A2(G132), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n835), .A2(G159), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1087), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1082), .B1(new_n1098), .B2(new_n818), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n913), .A2(new_n923), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n779), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n917), .A2(new_n922), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n654), .B(new_n812), .C1(new_n714), .C2(new_n717), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n861), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n871), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n914), .B(KEYINPUT114), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n708), .A2(G330), .A3(new_n931), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n915), .B1(new_n862), .B2(new_n871), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1110), .C1(new_n1101), .C2(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n930), .A2(G330), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n931), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1109), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1111), .B1(new_n913), .B2(new_n923), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1103), .B1(new_n1119), .B2(new_n1076), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT117), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n930), .A2(G330), .A3(new_n812), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n872), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1123), .A2(new_n861), .A3(new_n1105), .A4(new_n1110), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n708), .A2(G330), .A3(new_n812), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1125), .A2(new_n872), .B1(new_n1113), .B2(new_n931), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n1126), .B2(new_n863), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT116), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n462), .A2(new_n930), .A3(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT115), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n462), .A2(new_n930), .A3(KEYINPUT115), .A4(G330), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n927), .A2(new_n1128), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1131), .A2(new_n634), .A3(new_n926), .A4(new_n1132), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT116), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1127), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1119), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1112), .A2(new_n1118), .A3(new_n1136), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n676), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1120), .A2(KEYINPUT117), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1121), .A2(new_n1140), .A3(new_n1141), .ZN(G378));
  NAND2_X1  g0942(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n935), .A2(new_n929), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n939), .A2(new_n940), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(G330), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n633), .A2(new_n299), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n298), .A2(new_n653), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n925), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1146), .A2(new_n1147), .A3(G330), .A4(new_n1153), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1159));
  OAI211_X1 g0959(.A(KEYINPUT57), .B(new_n1145), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT121), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1145), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1153), .B1(new_n941), .B2(G330), .ZN(new_n1165));
  AND4_X1   g0965(.A1(G330), .A2(new_n1146), .A3(new_n1147), .A4(new_n1153), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n925), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT121), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT57), .A4(new_n1145), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1161), .A2(new_n1164), .A3(new_n676), .A4(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(G33), .A2(G41), .ZN(new_n1173));
  INV_X1    g0973(.A(G41), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G50), .B(new_n1173), .C1(new_n398), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(G128), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n757), .A2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n833), .A2(new_n749), .B1(new_n745), .B2(new_n1090), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G125), .C2(new_n740), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n1091), .B2(new_n756), .C1(new_n1004), .C2(new_n747), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g0981(.A(G124), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1173), .B1(new_n733), .B2(new_n1182), .C1(new_n840), .C2(new_n742), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1180), .B2(KEYINPUT59), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1175), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G41), .B(new_n255), .C1(new_n1041), .C2(G77), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n280), .B2(new_n742), .C1(new_n1031), .C2(new_n733), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT118), .Z(new_n1188));
  AOI22_X1  g0988(.A1(G116), .A2(new_n740), .B1(new_n828), .B2(G107), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n558), .B2(new_n749), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G68), .B2(new_n835), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(new_n1191), .C1(new_n319), .C2(new_n756), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT119), .Z(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1195));
  OAI21_X1  g0995(.A(new_n1185), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n818), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n727), .C1(G50), .C2(new_n820), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1154), .B2(new_n779), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1169), .B2(new_n726), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1172), .A2(new_n1202), .ZN(G375));
  INV_X1    g1003(.A(new_n1127), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1204), .A2(KEYINPUT122), .A3(new_n1076), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT122), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1127), .B2(new_n726), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n872), .A2(new_n779), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT123), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(KEYINPUT123), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n824), .A2(G116), .B1(G107), .B2(new_n764), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT124), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G283), .A2(new_n828), .B1(new_n734), .B2(G303), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n558), .B2(new_n745), .C1(new_n769), .C2(new_n739), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n398), .B1(new_n742), .B2(new_n257), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1212), .A2(new_n1044), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1058), .A2(new_n1090), .B1(new_n756), .B2(new_n1004), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n745), .A2(new_n840), .B1(new_n733), .B2(new_n1176), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n739), .A2(new_n833), .B1(new_n757), .B2(new_n1091), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n255), .B1(new_n747), .B2(new_n202), .C1(new_n280), .C2(new_n742), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n818), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n728), .C1(G68), .C2(new_n820), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT125), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1209), .A2(new_n1210), .A3(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1205), .A2(new_n1207), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n973), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1143), .A2(new_n1204), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1137), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(G381));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1172), .A2(new_n1231), .A3(new_n1202), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n988), .A2(new_n1012), .A3(new_n1080), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT126), .Z(new_n1235));
  OR4_X1    g1035(.A1(G381), .A2(new_n1232), .A3(new_n1233), .A4(new_n1235), .ZN(G407));
  INV_X1    g1036(.A(G343), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(G213), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT127), .Z(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(new_n1232), .C2(new_n1240), .ZN(G409));
  NAND3_X1  g1041(.A1(new_n1172), .A2(G378), .A3(new_n1202), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1202), .B1(new_n973), .B2(new_n1162), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1231), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1239), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1143), .A2(new_n1204), .A3(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n677), .B(new_n1136), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1226), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n848), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n848), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(G2897), .A3(new_n1239), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1239), .A2(G2897), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1253), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT63), .B1(new_n1245), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1254), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1245), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1245), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(new_n797), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1233), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1080), .B1(new_n988), .B2(new_n1012), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1266), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1264), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1233), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT61), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1262), .A2(new_n1263), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1245), .A2(new_n1274), .A3(new_n1260), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1245), .B2(new_n1258), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1274), .B1(new_n1245), .B2(new_n1260), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1275), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1271), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1273), .B1(new_n1279), .B2(new_n1280), .ZN(G405));
  XNOR2_X1  g1081(.A(new_n1271), .B(new_n1260), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G375), .B(new_n1231), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1282), .B(new_n1283), .ZN(G402));
endmodule


