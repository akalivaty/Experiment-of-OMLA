

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  NOR2_X2 U321 ( .A1(n425), .A2(n516), .ZN(n426) );
  INV_X1 U322 ( .A(G36GAT), .ZN(n350) );
  XNOR2_X1 U323 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U324 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U325 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n341) );
  XOR2_X1 U326 ( .A(n358), .B(n357), .Z(n565) );
  XOR2_X1 U327 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n289) );
  XOR2_X1 U328 ( .A(KEYINPUT27), .B(n457), .Z(n290) );
  XOR2_X1 U329 ( .A(G50GAT), .B(n342), .Z(n291) );
  INV_X1 U330 ( .A(KEYINPUT115), .ZN(n381) );
  XNOR2_X1 U331 ( .A(n381), .B(KEYINPUT47), .ZN(n382) );
  INV_X1 U332 ( .A(n396), .ZN(n317) );
  NOR2_X1 U333 ( .A1(n528), .A2(n458), .ZN(n459) );
  XNOR2_X1 U334 ( .A(n327), .B(KEYINPUT32), .ZN(n328) );
  XNOR2_X1 U335 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U336 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U337 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U338 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U339 ( .A(n336), .B(n335), .ZN(n340) );
  XNOR2_X1 U340 ( .A(n571), .B(n341), .ZN(n552) );
  XNOR2_X1 U341 ( .A(n326), .B(n325), .ZN(n575) );
  XOR2_X1 U342 ( .A(n443), .B(n442), .Z(n528) );
  XNOR2_X1 U343 ( .A(n490), .B(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U344 ( .A(n403), .B(n402), .ZN(n518) );
  XNOR2_X1 U345 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U346 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U347 ( .A(G197GAT), .B(KEYINPUT21), .Z(n392) );
  XOR2_X1 U348 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n293) );
  XNOR2_X1 U349 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n417) );
  XOR2_X1 U351 ( .A(n392), .B(n417), .Z(n295) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U353 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U354 ( .A(n296), .B(G211GAT), .Z(n300) );
  XOR2_X1 U355 ( .A(G162GAT), .B(KEYINPUT73), .Z(n298) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n368) );
  XNOR2_X1 U358 ( .A(n368), .B(KEYINPUT22), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U360 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n302) );
  XNOR2_X1 U361 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n301) );
  XNOR2_X1 U362 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U363 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U364 ( .A(G148GAT), .B(G204GAT), .Z(n306) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n329) );
  XNOR2_X1 U367 ( .A(G22GAT), .B(G155GAT), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n307), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n329), .B(n322), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n463) );
  XOR2_X1 U371 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n311) );
  XNOR2_X1 U372 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n310) );
  XNOR2_X1 U373 ( .A(n311), .B(n310), .ZN(n326) );
  XNOR2_X1 U374 ( .A(G71GAT), .B(G57GAT), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n312), .B(KEYINPUT13), .ZN(n338) );
  XOR2_X1 U376 ( .A(n338), .B(G64GAT), .Z(n314) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n314), .B(n313), .ZN(n320) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G1GAT), .ZN(n315) );
  XNOR2_X1 U380 ( .A(n315), .B(KEYINPUT67), .ZN(n342) );
  XNOR2_X1 U381 ( .A(n342), .B(G127GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .ZN(n316) );
  XNOR2_X1 U383 ( .A(n316), .B(G211GAT), .ZN(n396) );
  XOR2_X1 U384 ( .A(n321), .B(KEYINPUT14), .Z(n324) );
  XNOR2_X1 U385 ( .A(n322), .B(KEYINPUT79), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U387 ( .A(KEYINPUT113), .B(n575), .ZN(n560) );
  NAND2_X1 U388 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U389 ( .A(G99GAT), .B(G85GAT), .Z(n365) );
  XNOR2_X1 U390 ( .A(n330), .B(n365), .ZN(n336) );
  XOR2_X1 U391 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n332) );
  XNOR2_X1 U392 ( .A(KEYINPUT71), .B(KEYINPUT69), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n334) );
  XNOR2_X1 U394 ( .A(G120GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n337), .B(G64GAT), .ZN(n397) );
  XOR2_X1 U397 ( .A(n338), .B(n397), .Z(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n571) );
  INV_X1 U399 ( .A(n552), .ZN(n538) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n291), .B(n343), .ZN(n353) );
  XOR2_X1 U402 ( .A(G113GAT), .B(G141GAT), .Z(n345) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G197GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n347) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G8GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U409 ( .A(n354), .B(KEYINPUT66), .Z(n358) );
  XOR2_X1 U410 ( .A(G29GAT), .B(G43GAT), .Z(n356) );
  XNOR2_X1 U411 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n369) );
  XNOR2_X1 U413 ( .A(n369), .B(KEYINPUT68), .ZN(n357) );
  INV_X1 U414 ( .A(n565), .ZN(n535) );
  NAND2_X1 U415 ( .A1(n538), .A2(n535), .ZN(n360) );
  INV_X1 U416 ( .A(KEYINPUT46), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n361) );
  NOR2_X1 U418 ( .A1(n560), .A2(n361), .ZN(n362) );
  XNOR2_X1 U419 ( .A(KEYINPUT114), .B(n362), .ZN(n380) );
  XOR2_X1 U420 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n364) );
  XNOR2_X1 U421 ( .A(G134GAT), .B(KEYINPUT76), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n379) );
  XOR2_X1 U423 ( .A(KEYINPUT74), .B(n365), .Z(n367) );
  XOR2_X1 U424 ( .A(G36GAT), .B(G190GAT), .Z(n401) );
  XNOR2_X1 U425 ( .A(n401), .B(G92GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U428 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n371) );
  XNOR2_X1 U429 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n377) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U435 ( .A(n379), .B(n378), .Z(n545) );
  INV_X1 U436 ( .A(n545), .ZN(n558) );
  AND2_X1 U437 ( .A1(n380), .A2(n558), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U439 ( .A(KEYINPUT36), .B(n545), .Z(n579) );
  NOR2_X1 U440 ( .A1(n579), .A2(n575), .ZN(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT45), .B(n384), .Z(n385) );
  NOR2_X1 U442 ( .A1(n571), .A2(n385), .ZN(n386) );
  NAND2_X1 U443 ( .A1(n565), .A2(n386), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n389), .B(KEYINPUT48), .ZN(n530) );
  XNOR2_X1 U446 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n289), .B(n390), .ZN(n436) );
  XNOR2_X1 U448 ( .A(n436), .B(KEYINPUT91), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n391), .B(KEYINPUT90), .ZN(n395) );
  XNOR2_X1 U450 ( .A(G204GAT), .B(G218GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n395), .B(n394), .Z(n399) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U455 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  NAND2_X1 U457 ( .A1(n530), .A2(n518), .ZN(n405) );
  XOR2_X1 U458 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n425) );
  XOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT88), .Z(n407) );
  XNOR2_X1 U461 ( .A(KEYINPUT6), .B(KEYINPUT89), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n424) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G148GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U466 ( .A(KEYINPUT5), .B(G57GAT), .Z(n411) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(G155GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U469 ( .A(n413), .B(n412), .Z(n422) );
  XOR2_X1 U470 ( .A(G127GAT), .B(G134GAT), .Z(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U473 ( .A(G113GAT), .B(n416), .Z(n437) );
  XOR2_X1 U474 ( .A(n417), .B(KEYINPUT1), .Z(n419) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n437), .B(n420), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U479 ( .A(n424), .B(n423), .Z(n469) );
  INV_X1 U480 ( .A(n469), .ZN(n516) );
  XOR2_X1 U481 ( .A(KEYINPUT65), .B(n426), .Z(n564) );
  NAND2_X1 U482 ( .A1(n463), .A2(n564), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n427), .B(KEYINPUT55), .ZN(n444) );
  NAND2_X1 U484 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XOR2_X1 U485 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n429) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(KEYINPUT82), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U488 ( .A(G190GAT), .B(G99GAT), .Z(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n443) );
  XOR2_X1 U491 ( .A(G183GAT), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U494 ( .A(G71GAT), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n442) );
  AND2_X1 U498 ( .A1(n444), .A2(n528), .ZN(n561) );
  NAND2_X1 U499 ( .A1(n561), .A2(n538), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n446) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT56), .Z(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(G1349GAT) );
  NAND2_X1 U504 ( .A1(n561), .A2(n535), .ZN(n450) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(G1348GAT) );
  NAND2_X1 U507 ( .A1(n561), .A2(n545), .ZN(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n452) );
  INV_X1 U509 ( .A(G190GAT), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n476) );
  NOR2_X1 U511 ( .A1(n571), .A2(n565), .ZN(n455) );
  XOR2_X1 U512 ( .A(KEYINPUT72), .B(n455), .Z(n489) );
  NOR2_X1 U513 ( .A1(n545), .A2(n575), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT16), .ZN(n473) );
  XOR2_X1 U515 ( .A(n518), .B(KEYINPUT92), .Z(n457) );
  AND2_X1 U516 ( .A1(n516), .A2(n290), .ZN(n529) );
  XOR2_X1 U517 ( .A(n463), .B(KEYINPUT28), .Z(n523) );
  INV_X1 U518 ( .A(n523), .ZN(n532) );
  NAND2_X1 U519 ( .A1(n529), .A2(n532), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT93), .ZN(n472) );
  NAND2_X1 U521 ( .A1(n528), .A2(n518), .ZN(n460) );
  NAND2_X1 U522 ( .A1(n460), .A2(n463), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT95), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n463), .A2(n528), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(n563) );
  NAND2_X1 U528 ( .A1(n290), .A2(n563), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT96), .B(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n473), .A2(n486), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT97), .B(n474), .Z(n502) );
  NOR2_X1 U535 ( .A1(n489), .A2(n502), .ZN(n484) );
  NAND2_X1 U536 ( .A1(n484), .A2(n516), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U538 ( .A(G1GAT), .B(n477), .Z(G1324GAT) );
  XOR2_X1 U539 ( .A(G8GAT), .B(KEYINPUT99), .Z(n479) );
  NAND2_X1 U540 ( .A1(n484), .A2(n518), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n481) );
  NAND2_X1 U543 ( .A1(n484), .A2(n528), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(n483) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT100), .Z(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n484), .A2(n523), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n492) );
  NAND2_X1 U550 ( .A1(n486), .A2(n575), .ZN(n487) );
  NOR2_X1 U551 ( .A1(n579), .A2(n487), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n488), .B(KEYINPUT37), .ZN(n515) );
  NOR2_X1 U553 ( .A1(n515), .A2(n489), .ZN(n490) );
  NAND2_X1 U554 ( .A1(n499), .A2(n516), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  XOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT103), .Z(n495) );
  NAND2_X1 U558 ( .A1(n518), .A2(n499), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U561 ( .A1(n499), .A2(n528), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U563 ( .A(n498), .B(G43GAT), .Z(G1330GAT) );
  XOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT105), .Z(n501) );
  NAND2_X1 U565 ( .A1(n523), .A2(n499), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NAND2_X1 U568 ( .A1(n565), .A2(n538), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n502), .A2(n514), .ZN(n509) );
  NAND2_X1 U570 ( .A1(n509), .A2(n516), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n518), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U575 ( .A1(n509), .A2(n528), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U579 ( .A1(n509), .A2(n523), .ZN(n510) );
  XNOR2_X1 U580 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT109), .Z(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n524), .A2(n516), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  XOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT111), .Z(n522) );
  NAND2_X1 U590 ( .A1(n524), .A2(n528), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n522), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n526) );
  NAND2_X1 U593 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT117), .Z(n537) );
  INV_X1 U597 ( .A(n528), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n531), .Z(n550) );
  NAND2_X1 U600 ( .A1(n550), .A2(n532), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U605 ( .A1(n546), .A2(n538), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n542) );
  NAND2_X1 U609 ( .A1(n546), .A2(n560), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n563), .A2(n550), .ZN(n557) );
  NOR2_X1 U617 ( .A1(n565), .A2(n557), .ZN(n551) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n557), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G148GAT), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n575), .A2(n557), .ZN(n556) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n559), .Z(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n578) );
  NOR2_X1 U630 ( .A1(n565), .A2(n578), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT125), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U637 ( .A(n578), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

