//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n455), .A2(new_n459), .B1(new_n450), .B2(new_n456), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n462), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G101), .A3(G2104), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  AND3_X1   g056(.A1(new_n469), .A2(new_n478), .A3(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n477), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n462), .A2(G138), .A3(new_n479), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n472), .B2(new_n474), .ZN(new_n493));
  AND2_X1   g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n475), .A2(KEYINPUT4), .A3(G138), .ZN(new_n497));
  NAND2_X1  g072(.A1(G102), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n496), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(G62), .A3(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT72), .A3(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT71), .B1(new_n511), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n513), .A2(new_n517), .A3(new_n506), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n507), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n517), .A2(new_n510), .A3(new_n512), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n501), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(G166));
  AND3_X1   g101(.A1(new_n513), .A2(G543), .A3(new_n517), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT74), .B(G89), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n518), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n509), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n527), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n509), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n518), .A2(G81), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT75), .B(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n527), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  AND3_X1   g130(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT77), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT77), .B1(new_n502), .B2(new_n504), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT76), .Z(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n522), .A2(G91), .A3(new_n506), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n522), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n517), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n567), .ZN(G299));
  INV_X1    g143(.A(G166), .ZN(G303));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n519), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n506), .A2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n527), .A2(G49), .B1(new_n573), .B2(G651), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n518), .A2(KEYINPUT78), .A3(G87), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n527), .A2(G48), .B1(new_n518), .B2(G86), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n505), .A2(KEYINPUT79), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n505), .B2(new_n578), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n527), .A2(G47), .B1(new_n518), .B2(G85), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT80), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n509), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n518), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n556), .A2(new_n557), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G66), .ZN(new_n595));
  INV_X1    g170(.A(G79), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n501), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NOR2_X1   g183(.A1(new_n549), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n600), .A2(new_n607), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n483), .A2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n477), .A2(G135), .ZN(new_n615));
  NOR2_X1   g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(new_n479), .B2(G111), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  XOR2_X1   g194(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n620));
  NOR3_X1   g195(.A1(new_n470), .A2(new_n471), .A3(G2105), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT13), .B(G2100), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT84), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2451), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G14), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT85), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2072), .B(G2078), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT86), .Z(new_n648));
  XOR2_X1   g223(.A(new_n646), .B(KEYINPUT17), .Z(new_n649));
  INV_X1    g224(.A(new_n645), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n649), .A3(new_n642), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n642), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT87), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G21), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G168), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1966), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT31), .B(G11), .Z(new_n683));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(G28), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(G28), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n618), .A2(new_n687), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT95), .Z(new_n691));
  INV_X1    g266(.A(G1961), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT96), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G5), .B2(G16), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n693), .A2(G5), .A3(G16), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n694), .B(new_n695), .C1(G301), .C2(new_n679), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n689), .B(new_n691), .C1(new_n692), .C2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT97), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G160), .A2(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(KEYINPUT24), .A2(G34), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  AOI21_X1  g278(.A(G29), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT93), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT93), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT94), .B(G2084), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n483), .ZN(new_n710));
  INV_X1    g285(.A(G128), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n710), .A2(KEYINPUT91), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(new_n479), .B2(G116), .ZN(new_n713));
  INV_X1    g288(.A(G104), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n479), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n477), .B2(G140), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT91), .B1(new_n710), .B2(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n687), .A2(G26), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2067), .ZN(new_n724));
  INV_X1    g299(.A(G2078), .ZN(new_n725));
  NAND2_X1  g300(.A1(G164), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G27), .B2(G29), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n679), .A2(KEYINPUT23), .A3(G20), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT23), .ZN(new_n730));
  INV_X1    g305(.A(G20), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n732), .C1(new_n604), .C2(new_n679), .ZN(new_n733));
  INV_X1    g308(.A(G1956), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n699), .A2(new_n709), .A3(new_n728), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n687), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n687), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2090), .ZN(new_n740));
  INV_X1    g315(.A(G1341), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n549), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G16), .B2(G19), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n740), .B1(new_n741), .B2(new_n743), .C1(new_n725), .C2(new_n727), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n477), .A2(G139), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  AOI22_X1  g322(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n747), .C1(new_n479), .C2(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G33), .B(new_n749), .S(G29), .Z(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2072), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n696), .A2(new_n692), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n707), .A2(new_n708), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n736), .A2(new_n744), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n687), .A2(G32), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n477), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n483), .A2(G129), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n479), .A2(G105), .A3(G2104), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND4_X1  g336(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(new_n687), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n743), .A2(new_n741), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G23), .ZN(new_n768));
  INV_X1    g343(.A(G288), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT33), .B(G1976), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G6), .B(G305), .S(G16), .Z(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT32), .B(G1981), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT90), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n679), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n679), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n772), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT34), .Z(new_n782));
  AOI22_X1  g357(.A1(G119), .A2(new_n483), .B1(new_n477), .B2(G131), .ZN(new_n783));
  OR2_X1    g358(.A1(G95), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT88), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G25), .B(new_n787), .S(G29), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT35), .B(G1991), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT89), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G290), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(new_n679), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n679), .B2(G24), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n782), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT36), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n755), .A2(new_n766), .A3(new_n767), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n679), .A2(G4), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n600), .B2(new_n679), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1348), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n800), .A2(KEYINPUT98), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT98), .B1(new_n800), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n800), .A2(new_n807), .A3(new_n803), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n800), .B2(new_n803), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(G150));
  NAND2_X1  g385(.A1(new_n518), .A2(G93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n527), .A2(G55), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n811), .B(new_n812), .C1(new_n509), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  XOR2_X1   g391(.A(new_n814), .B(new_n548), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n599), .A2(new_n607), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(G860), .ZN(G145));
  XNOR2_X1  g397(.A(new_n718), .B(G164), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G160), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n488), .B(KEYINPUT100), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n618), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n749), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n483), .A2(G130), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n477), .A2(G142), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n479), .A2(G118), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT101), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n762), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n787), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n622), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n828), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT102), .B(G37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g416(.A(new_n599), .B(G299), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT41), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n610), .B(new_n817), .ZN(new_n844));
  MUX2_X1   g419(.A(new_n842), .B(new_n843), .S(new_n844), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT42), .ZN(new_n846));
  XNOR2_X1  g421(.A(G288), .B(G166), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G290), .ZN(new_n848));
  XNOR2_X1  g423(.A(G305), .B(KEYINPUT103), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n846), .B(new_n850), .Z(new_n851));
  MUX2_X1   g426(.A(new_n814), .B(new_n851), .S(G868), .Z(G295));
  MUX2_X1   g427(.A(new_n814), .B(new_n851), .S(G868), .Z(G331));
  XOR2_X1   g428(.A(G286), .B(G301), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n817), .B(new_n854), .ZN(new_n855));
  MUX2_X1   g430(.A(new_n842), .B(new_n843), .S(new_n855), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n850), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(KEYINPUT43), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n839), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT44), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n859), .A2(new_n862), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n861), .A2(KEYINPUT43), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g443(.A(KEYINPUT126), .ZN(new_n869));
  INV_X1    g444(.A(G1384), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n496), .B2(new_n499), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT104), .B(G40), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n469), .A2(new_n478), .A3(new_n481), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(G1996), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n763), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT105), .ZN(new_n880));
  INV_X1    g455(.A(G2067), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n718), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G1996), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n763), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n880), .B1(new_n876), .B2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n787), .B(new_n789), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT106), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n877), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n792), .A2(new_n795), .ZN(new_n889));
  NAND2_X1  g464(.A1(G290), .A2(G1986), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n877), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n875), .A2(new_n871), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(G8), .ZN(new_n896));
  OAI21_X1  g471(.A(G8), .B1(new_n875), .B2(new_n871), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT110), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT49), .ZN(new_n900));
  NOR2_X1   g475(.A1(G305), .A2(G1981), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G1981), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n577), .B2(new_n583), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n900), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n901), .A2(KEYINPUT49), .A3(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT52), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n896), .A2(new_n898), .B1(G1976), .B2(new_n769), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G1976), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT52), .B1(G288), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n875), .ZN(new_n916));
  OAI211_X1 g491(.A(KEYINPUT45), .B(new_n870), .C1(new_n496), .C2(new_n499), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n873), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT107), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(new_n873), .A3(new_n920), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n779), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT50), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n871), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT50), .B(new_n870), .C1(new_n496), .C2(new_n499), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n916), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(G2090), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(KEYINPUT108), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  AOI21_X1  g507(.A(G1971), .B1(new_n919), .B2(new_n921), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(G8), .ZN(new_n935));
  NOR2_X1   g510(.A1(G166), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(G166), .B2(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n931), .A2(new_n934), .A3(G8), .A4(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n915), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(G8), .B1(new_n933), .B2(new_n929), .ZN(new_n944));
  INV_X1    g519(.A(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n922), .B2(G2078), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n916), .A2(new_n873), .A3(new_n917), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(KEYINPUT53), .A3(new_n725), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n928), .A2(KEYINPUT115), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n875), .B1(new_n925), .B2(new_n926), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT115), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(KEYINPUT122), .B(G1961), .Z(new_n956));
  NAND3_X1  g531(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n949), .A2(new_n951), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT62), .ZN(new_n960));
  INV_X1    g535(.A(G2084), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n927), .A2(new_n961), .A3(new_n916), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n963));
  INV_X1    g538(.A(G1966), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n918), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n953), .A2(new_n966), .A3(new_n961), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n963), .A2(G168), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G8), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G8), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n972), .B2(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(G286), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n969), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n971), .B2(G8), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n976), .A2(new_n978), .A3(new_n970), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n960), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n969), .ZN(new_n981));
  INV_X1    g556(.A(new_n974), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n982), .A2(new_n978), .A3(new_n970), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT62), .B(new_n981), .C1(new_n983), .C2(new_n969), .ZN(new_n984));
  AOI211_X1 g559(.A(G301), .B(new_n959), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n561), .B1(new_n594), .B2(G65), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n563), .B1(new_n987), .B2(new_n509), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n564), .A2(new_n567), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT114), .ZN(new_n991));
  NOR2_X1   g566(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  NAND3_X1  g568(.A1(G299), .A2(new_n993), .A3(new_n986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(new_n994), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n993), .B1(G299), .B2(new_n986), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n953), .A2(G1956), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT56), .B(G2072), .ZN(new_n1001));
  AND4_X1   g576(.A1(new_n873), .A2(new_n916), .A3(new_n917), .A4(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n995), .B(new_n999), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1348), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n952), .A2(new_n1004), .A3(new_n955), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n894), .A2(G2067), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n928), .A2(new_n734), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n950), .A2(new_n1001), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n997), .A2(new_n998), .A3(new_n996), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1011), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1010), .A2(new_n600), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(KEYINPUT61), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1003), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n916), .A2(new_n873), .A3(new_n883), .A4(new_n917), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT58), .B(G1341), .Z(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n875), .B2(new_n871), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1023), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n549), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT118), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(KEYINPUT118), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n549), .B(new_n1032), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1015), .A2(new_n1003), .A3(new_n1017), .A4(KEYINPUT61), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1021), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1028), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n548), .B1(new_n1039), .B2(new_n1026), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1033), .A2(new_n1031), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n1021), .A4(new_n1036), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1008), .A2(new_n1009), .A3(KEYINPUT60), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT60), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n600), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT60), .B(new_n599), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1003), .B(new_n1016), .C1(new_n1046), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n949), .A2(new_n957), .ZN(new_n1053));
  XNOR2_X1  g628(.A(G301), .B(KEYINPUT54), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n725), .A2(KEYINPUT53), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n873), .A2(G40), .A3(G160), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(KEYINPUT124), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n917), .C1(KEYINPUT124), .C2(new_n1057), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1055), .A2(new_n1059), .B1(new_n1054), .B2(new_n958), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n943), .A2(new_n1060), .A3(new_n946), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n975), .A2(new_n979), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n947), .A2(new_n985), .B1(new_n1052), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n972), .A2(G286), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n931), .A2(G8), .A3(new_n934), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n945), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n943), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n915), .A2(new_n942), .A3(new_n946), .A4(new_n1066), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1067), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n908), .A2(new_n912), .A3(new_n769), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n902), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n899), .ZN(new_n1076));
  INV_X1    g651(.A(new_n915), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n942), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1065), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT112), .B(new_n1078), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n893), .B1(new_n1064), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n889), .A2(new_n877), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT125), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT48), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n888), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n787), .A2(new_n789), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n885), .A2(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n718), .A2(G2067), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n877), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n878), .A2(KEYINPUT46), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n878), .A2(KEYINPUT46), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n882), .A2(new_n763), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1092), .B(new_n1093), .C1(new_n877), .C2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1095), .B(KEYINPUT47), .Z(new_n1096));
  NOR3_X1   g671(.A1(new_n1087), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n869), .B1(new_n1083), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1052), .A2(new_n1063), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT112), .ZN(new_n1102));
  AOI21_X1  g677(.A(G301), .B1(new_n980), .B2(new_n984), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n947), .A3(new_n958), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1073), .A2(new_n1065), .A3(new_n1079), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n892), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT126), .A3(new_n1097), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1099), .A2(new_n1108), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g684(.A1(new_n865), .A2(new_n866), .ZN(new_n1111));
  OR4_X1    g685(.A1(new_n460), .A2(G401), .A3(G227), .A4(G229), .ZN(new_n1112));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n1113));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g688(.A(new_n1114), .B1(new_n839), .B2(new_n838), .ZN(new_n1115));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1116));
  AND3_X1   g690(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .ZN(G308));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .ZN(G225));
endmodule


