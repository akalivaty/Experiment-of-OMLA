//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  AND2_X1   g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT70), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(KEYINPUT70), .A3(new_n464), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(new_n470), .B1(G113), .B2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(KEYINPUT69), .B(G125), .C1(new_n461), .C2(new_n462), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n461), .A2(new_n462), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n460), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n477), .B(new_n481), .C1(G124), .C2(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n485));
  INV_X1    g060(.A(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n460), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n495), .B(new_n496), .C1(new_n462), .C2(new_n461), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n496), .B1(new_n499), .B2(new_n495), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n493), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n495), .B1(new_n461), .B2(new_n462), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n497), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n493), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT73), .Z(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n509), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  AND2_X1   g101(.A1(new_n517), .A2(new_n520), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n529), .B(new_n531), .C1(new_n532), .C2(new_n523), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(new_n517), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  INV_X1    g111(.A(G77), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n512), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n540), .B1(new_n537), .B2(new_n512), .C1(new_n535), .C2(new_n536), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(G651), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n520), .A2(G543), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n527), .A2(G90), .B1(new_n543), .B2(G52), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n509), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n527), .A2(G81), .B1(new_n543), .B2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT75), .Z(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND3_X1  g131(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n509), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n527), .A2(G91), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(new_n542), .A2(new_n544), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n543), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n517), .A2(G87), .A3(new_n520), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n509), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n521), .A2(new_n572), .B1(new_n523), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n509), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n527), .A2(G85), .B1(new_n543), .B2(G47), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G79), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G66), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n535), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G54), .B2(new_n543), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n517), .A2(G92), .A3(new_n520), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G171), .B2(new_n589), .ZN(G284));
  OAI21_X1  g166(.A(new_n590), .B1(G171), .B2(new_n589), .ZN(G321));
  NAND2_X1  g167(.A1(G299), .A2(new_n589), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n589), .B2(G168), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(new_n589), .B2(G168), .ZN(G280));
  INV_X1    g170(.A(new_n588), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT76), .B(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(G860), .B2(new_n597), .ZN(G148));
  NOR2_X1   g173(.A1(new_n550), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n597), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT77), .Z(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g178(.A1(new_n482), .A2(G123), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT80), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n479), .A2(G135), .ZN(new_n606));
  NOR3_X1   g181(.A1(new_n460), .A2(KEYINPUT81), .A3(G111), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT81), .B1(new_n460), .B2(G111), .ZN(new_n608));
  OR2_X1    g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n608), .A2(G2104), .A3(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n610), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(G2096), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n485), .A2(new_n486), .A3(G2105), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT79), .B(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n611), .A2(G2096), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n612), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT83), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n628), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n640), .ZN(new_n647));
  INV_X1    g222(.A(new_n641), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n643), .A3(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(new_n642), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n657), .A2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n665));
  OAI221_X1 g240(.A(new_n663), .B1(new_n657), .B2(new_n662), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n664), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1981), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  NAND2_X1  g248(.A1(G288), .A2(KEYINPUT89), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n675));
  NAND4_X1  g250(.A1(new_n566), .A2(new_n675), .A3(new_n567), .A4(new_n568), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G16), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G16), .B2(G23), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT87), .B(G16), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n575), .B2(G16), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n682), .A2(new_n683), .A3(new_n689), .A4(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n695));
  MUX2_X1   g270(.A(G24), .B(G290), .S(new_n685), .Z(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT88), .Z(new_n697));
  INV_X1    g272(.A(G1986), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n479), .A2(G131), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n482), .A2(G119), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n460), .A2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT86), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n699), .A2(new_n700), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n695), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT36), .ZN(new_n713));
  NOR2_X1   g288(.A1(G4), .A2(G16), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n588), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1348), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n685), .A2(G19), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n550), .B2(new_n685), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1341), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G26), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n479), .A2(G140), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n482), .A2(G128), .ZN(new_n727));
  OR2_X1    g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n723), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n719), .A2(new_n722), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  NOR2_X1   g310(.A1(G27), .A2(G29), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G164), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2078), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n684), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NOR2_X1   g318(.A1(G5), .A2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G301), .B2(new_n716), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n742), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n738), .B(new_n747), .C1(new_n743), .C2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n723), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n723), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT29), .Z(new_n751));
  INV_X1    g326(.A(G2090), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n723), .B1(KEYINPUT24), .B2(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(KEYINPUT24), .B2(G34), .ZN(new_n756));
  INV_X1    g331(.A(G160), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n753), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(G29), .A2(G33), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n479), .A2(G139), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT92), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n460), .C2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(new_n723), .ZN(new_n767));
  INV_X1    g342(.A(G2072), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n479), .A2(G141), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT26), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n772), .B(new_n774), .C1(G129), .C2(new_n482), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n723), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n723), .B2(G32), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n769), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n758), .A2(new_n754), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n751), .B2(new_n752), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT31), .B(G11), .Z(new_n785));
  NOR2_X1   g360(.A1(new_n611), .A2(new_n723), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT30), .B(G28), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n785), .B(new_n786), .C1(new_n723), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n716), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n767), .A2(new_n768), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n759), .A2(new_n782), .A3(new_n784), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n713), .A2(new_n735), .A3(new_n748), .A4(new_n795), .ZN(G150));
  INV_X1    g371(.A(G150), .ZN(G311));
  AOI22_X1  g372(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(new_n509), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n527), .A2(G93), .B1(new_n543), .B2(G55), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G860), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n799), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n805), .B1(new_n799), .B2(new_n800), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n807), .A2(new_n549), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n550), .B1(new_n810), .B2(new_n806), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G559), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT96), .B1(new_n588), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT38), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(KEYINPUT38), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n820), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n822), .A2(new_n812), .A3(new_n818), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT98), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n824), .A2(new_n830), .A3(new_n825), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n827), .A2(KEYINPUT99), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT99), .B1(new_n827), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n804), .B1(new_n833), .B2(new_n834), .ZN(G145));
  NAND2_X1  g410(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n776), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n705), .B(new_n615), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n840), .B1(new_n490), .B2(new_n491), .C1(new_n478), .C2(new_n484), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT103), .B1(new_n489), .B2(new_n492), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n506), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n730), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n482), .A2(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n460), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n479), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n839), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n611), .B(G162), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n757), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(G37), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n851), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g433(.A(new_n549), .B1(new_n807), .B2(new_n808), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n810), .A2(new_n550), .A3(new_n806), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n600), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n600), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n560), .A2(new_n561), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n588), .A2(new_n558), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n585), .B(KEYINPUT10), .ZN(new_n867));
  NAND3_X1  g442(.A1(G299), .A2(new_n867), .A3(new_n584), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n596), .A2(KEYINPUT105), .A3(G299), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT41), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n865), .A2(new_n872), .A3(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT106), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT106), .B1(new_n869), .B2(new_n870), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n879));
  NAND3_X1  g454(.A1(G303), .A2(new_n578), .A3(new_n579), .ZN(new_n880));
  NAND2_X1  g455(.A1(G290), .A2(G166), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n677), .A2(new_n575), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n677), .A2(new_n575), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n678), .A2(G305), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n887), .A2(new_n881), .A3(new_n880), .A4(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n879), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(KEYINPUT108), .B(new_n890), .C1(new_n886), .C2(new_n888), .ZN(new_n893));
  OAI221_X1 g468(.A(new_n875), .B1(new_n878), .B2(new_n863), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n875), .B1(new_n878), .B2(new_n863), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n894), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n801), .A2(new_n589), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n901), .A2(new_n904), .A3(new_n902), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  INV_X1    g483(.A(new_n874), .ZN(new_n909));
  NAND2_X1  g484(.A1(G301), .A2(G286), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(G301), .A2(G286), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n860), .B(new_n859), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G171), .A2(G168), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n910), .B(new_n914), .C1(new_n809), .C2(new_n811), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT110), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n910), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n812), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n909), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n913), .A2(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n869), .A2(new_n870), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n889), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n917), .ZN(new_n927));
  INV_X1    g502(.A(new_n919), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n878), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n865), .A2(new_n868), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n922), .A2(new_n872), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n921), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n921), .A2(new_n932), .A3(KEYINPUT111), .A4(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n889), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n908), .B1(new_n940), .B2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n924), .A2(new_n925), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n889), .B1(new_n920), .B2(new_n923), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n926), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n942), .B2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT112), .B1(new_n949), .B2(new_n908), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n951), .B(KEYINPUT44), .C1(new_n947), .C2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n950), .B2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n843), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n463), .A2(KEYINPUT70), .A3(new_n464), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(new_n465), .ZN(new_n959));
  NAND2_X1  g534(.A1(G113), .A2(G2104), .ZN(new_n960));
  INV_X1    g535(.A(G125), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n487), .B2(new_n488), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n962), .B2(KEYINPUT69), .ZN(new_n963));
  INV_X1    g538(.A(new_n472), .ZN(new_n964));
  OAI21_X1  g539(.A(G2105), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n959), .A2(new_n965), .A3(G40), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n968), .A2(G1986), .A3(G290), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT48), .Z(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n776), .B(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n730), .B(G2067), .Z(new_n973));
  INV_X1    g548(.A(new_n708), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n705), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n705), .A2(new_n974), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n972), .A2(new_n973), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n970), .B1(new_n978), .B2(new_n968), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n973), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n980), .A2(new_n975), .B1(G2067), .B2(new_n730), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n967), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n967), .A2(new_n971), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n777), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n967), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n985), .B2(new_n984), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n979), .B(new_n982), .C1(new_n983), .C2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n983), .B2(new_n988), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n503), .A2(new_n954), .A3(new_n507), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n956), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n468), .A2(new_n473), .A3(new_n994), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n478), .A2(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n996));
  AOI22_X1  g571(.A1(KEYINPUT103), .A2(new_n996), .B1(new_n505), .B2(new_n497), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n997), .B2(new_n841), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n991), .B1(new_n1000), .B2(G2078), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n954), .A4(new_n507), .ZN(new_n1003));
  INV_X1    g578(.A(G2078), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n957), .A2(new_n1003), .A3(new_n995), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT125), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n843), .B2(new_n954), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(new_n966), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT125), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n1004), .A4(new_n1003), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(KEYINPUT53), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n966), .B1(new_n1012), .B2(new_n998), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n743), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT126), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT126), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1002), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n674), .A2(G1976), .A3(new_n676), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(G8), .C1(new_n966), .C2(new_n955), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT52), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n966), .A2(new_n955), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n575), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(G1981), .B1(new_n571), .B2(new_n574), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1032), .B(new_n1033), .C1(new_n1034), .C2(KEYINPUT49), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1033), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n571), .A2(new_n574), .A3(G1981), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1027), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1024), .A2(new_n1030), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n956), .B2(new_n992), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1971), .B1(new_n1043), .B2(new_n995), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n503), .A2(new_n1012), .A3(new_n954), .A4(new_n507), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n995), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G2090), .ZN(new_n1048));
  OAI21_X1  g623(.A(G8), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1050), .B2(KEYINPUT55), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G166), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(KEYINPUT55), .ZN(new_n1053));
  XOR2_X1   g628(.A(new_n1053), .B(KEYINPUT115), .Z(new_n1054));
  XOR2_X1   g629(.A(new_n1052), .B(new_n1054), .Z(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1041), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1013), .A2(new_n752), .A3(new_n1014), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1044), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1000), .A2(new_n688), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1013), .A2(new_n752), .A3(new_n1014), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT113), .A3(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(G8), .A3(new_n1055), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1021), .A2(new_n1065), .A3(G301), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n957), .A2(new_n1003), .A3(new_n995), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n791), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT117), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1070), .A3(new_n791), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1013), .A2(new_n754), .A3(new_n1014), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G286), .A2(G8), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT124), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1073), .B2(G8), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(KEYINPUT51), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1079), .B(new_n1075), .C1(new_n1073), .C2(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT62), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n754), .A2(new_n1082), .B1(new_n1068), .B2(KEYINPUT117), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1026), .B1(new_n1083), .B2(new_n1071), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1084), .B2(new_n1075), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1077), .A2(KEYINPUT51), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1076), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1066), .A2(new_n1081), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1041), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1064), .A2(new_n1084), .A3(G168), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1026), .B1(new_n1094), .B2(new_n1058), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1055), .B1(new_n1095), .B2(new_n1063), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1090), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1966), .B1(new_n1008), .B2(new_n1003), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1072), .B1(new_n1098), .B2(new_n1070), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1071), .ZN(new_n1100));
  OAI211_X1 g675(.A(G8), .B(G168), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1101), .A2(new_n1091), .A3(new_n1041), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1060), .A2(G8), .A3(new_n1063), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1056), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n1104), .A4(new_n1064), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1091), .B1(new_n1065), .B2(new_n1101), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1064), .A2(new_n1041), .ZN(new_n1108));
  INV_X1    g683(.A(G288), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1040), .A2(new_n1028), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1032), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1027), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1089), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1042), .A2(new_n1007), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n1116));
  NOR4_X1   g691(.A1(new_n473), .A2(new_n991), .A3(new_n994), .A4(G2078), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1016), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1001), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G171), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1001), .A2(G301), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT54), .B(new_n1121), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1085), .A2(new_n1086), .A3(new_n1076), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1064), .A4(new_n1057), .ZN(new_n1126));
  OAI21_X1  g701(.A(G171), .B1(new_n1122), .B2(new_n1002), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(G301), .A3(new_n1001), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT54), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  INV_X1    g706(.A(G1956), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1047), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n993), .A2(new_n995), .A3(new_n999), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G299), .B(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n966), .A2(new_n955), .A3(G2067), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1015), .B2(new_n718), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n588), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .A4(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n966), .A2(G1996), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n993), .A2(new_n999), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n995), .A2(new_n998), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n549), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1043), .A2(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT121), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(G1348), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n596), .A4(new_n1141), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n588), .B1(new_n1142), .B2(KEYINPUT60), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1163), .B2(new_n1141), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1140), .A2(KEYINPUT61), .A3(new_n1144), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1157), .A2(new_n1159), .A3(KEYINPUT122), .A4(KEYINPUT59), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1162), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT61), .B1(new_n1148), .B2(new_n1140), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1131), .B(new_n1149), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1148), .A2(new_n1140), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1141), .ZN(new_n1178));
  OAI211_X1 g753(.A(KEYINPUT60), .B(new_n1178), .C1(new_n1082), .C2(G1348), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(new_n1167), .A3(new_n596), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1165), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1169), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1151), .A2(KEYINPUT121), .A3(new_n1154), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT121), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1184));
  NAND2_X1  g759(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1185));
  NOR4_X1   g760(.A1(new_n1183), .A2(new_n1184), .A3(new_n549), .A4(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1161), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1177), .A2(new_n1182), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1131), .B1(new_n1190), .B2(new_n1149), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1174), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1113), .B1(new_n1130), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G290), .B(new_n698), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n968), .B1(new_n978), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n990), .B1(new_n1193), .B2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(new_n458), .ZN(new_n1198));
  NOR4_X1   g772(.A1(G229), .A2(new_n1198), .A3(G401), .A4(G227), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n1199), .A2(new_n857), .A3(new_n949), .ZN(G225));
  INV_X1    g774(.A(G225), .ZN(G308));
endmodule


