

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721;

  NOR2_X1 U367 ( .A1(n567), .A2(n566), .ZN(n593) );
  OR2_X2 U368 ( .A1(n565), .A2(n531), .ZN(n518) );
  BUF_X1 U369 ( .A(G953), .Z(n343) );
  XNOR2_X1 U370 ( .A(n480), .B(KEYINPUT72), .ZN(n452) );
  XNOR2_X1 U371 ( .A(n404), .B(n427), .ZN(n469) );
  AND2_X2 U372 ( .A1(n397), .A2(n395), .ZN(n548) );
  XNOR2_X1 U373 ( .A(n470), .B(n471), .ZN(n685) );
  AND2_X2 U374 ( .A1(n623), .A2(n622), .ZN(n625) );
  NOR2_X2 U375 ( .A1(n518), .A2(n571), .ZN(n559) );
  BUF_X1 U376 ( .A(G146), .Z(n355) );
  OR2_X2 U377 ( .A1(n672), .A2(G902), .ZN(n391) );
  XNOR2_X2 U378 ( .A(n435), .B(KEYINPUT3), .ZN(n482) );
  XNOR2_X2 U379 ( .A(G119), .B(G116), .ZN(n435) );
  XNOR2_X2 U380 ( .A(n441), .B(n392), .ZN(n451) );
  XNOR2_X2 U381 ( .A(n487), .B(n486), .ZN(n555) );
  XNOR2_X2 U382 ( .A(n708), .B(G101), .ZN(n480) );
  NOR2_X1 U383 ( .A1(n503), .A2(n530), .ZN(n360) );
  AND2_X1 U384 ( .A1(n376), .A2(n670), .ZN(n375) );
  XNOR2_X1 U385 ( .A(n368), .B(n367), .ZN(n580) );
  INV_X1 U386 ( .A(KEYINPUT35), .ZN(n387) );
  NOR2_X2 U387 ( .A1(n718), .A2(n719), .ZN(n578) );
  AND2_X1 U388 ( .A1(n720), .A2(n654), .ZN(n397) );
  XNOR2_X1 U389 ( .A(n388), .B(n387), .ZN(n720) );
  NAND2_X1 U390 ( .A1(n389), .A2(n587), .ZN(n388) );
  NOR2_X2 U391 ( .A1(n581), .A2(n580), .ZN(n660) );
  XNOR2_X1 U392 ( .A(n672), .B(n675), .ZN(n676) );
  XNOR2_X1 U393 ( .A(n432), .B(G478), .ZN(n544) );
  XNOR2_X1 U394 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n427) );
  NAND2_X1 U395 ( .A1(n710), .A2(G234), .ZN(n404) );
  INV_X4 U396 ( .A(G953), .ZN(n699) );
  XNOR2_X1 U397 ( .A(G125), .B(KEYINPUT10), .ZN(n462) );
  XOR2_X1 U398 ( .A(n424), .B(n423), .Z(n543) );
  NOR2_X1 U399 ( .A1(n633), .A2(G902), .ZN(n424) );
  INV_X1 U400 ( .A(G469), .ZN(n390) );
  INV_X1 U401 ( .A(n607), .ZN(n359) );
  AND2_X1 U402 ( .A1(n533), .A2(KEYINPUT22), .ZN(n402) );
  NOR2_X1 U403 ( .A1(G237), .A2(G902), .ZN(n446) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n382) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n353) );
  INV_X1 U406 ( .A(G134), .ZN(n392) );
  XNOR2_X1 U407 ( .A(n441), .B(n693), .ZN(n442) );
  XNOR2_X1 U408 ( .A(n385), .B(n384), .ZN(n439) );
  XNOR2_X1 U409 ( .A(KEYINPUT17), .B(KEYINPUT90), .ZN(n384) );
  XNOR2_X1 U410 ( .A(n592), .B(n383), .ZN(n561) );
  INV_X1 U411 ( .A(KEYINPUT38), .ZN(n383) );
  XNOR2_X1 U412 ( .A(n420), .B(n419), .ZN(n633) );
  XNOR2_X1 U413 ( .A(n363), .B(n413), .ZN(n420) );
  NAND2_X1 U414 ( .A1(n488), .A2(n599), .ZN(n361) );
  NOR2_X1 U415 ( .A1(n370), .A2(n359), .ZN(n358) );
  NOR2_X1 U416 ( .A1(n655), .A2(n659), .ZN(n586) );
  XNOR2_X1 U417 ( .A(n576), .B(KEYINPUT46), .ZN(n577) );
  XNOR2_X1 U418 ( .A(n386), .B(KEYINPUT93), .ZN(n385) );
  XNOR2_X1 U419 ( .A(KEYINPUT78), .B(G125), .ZN(n386) );
  NAND2_X1 U420 ( .A1(G234), .A2(G237), .ZN(n490) );
  NAND2_X1 U421 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U422 ( .A(KEYINPUT87), .ZN(n377) );
  INV_X1 U423 ( .A(n671), .ZN(n378) );
  AND2_X1 U424 ( .A1(n671), .A2(KEYINPUT87), .ZN(n380) );
  XNOR2_X1 U425 ( .A(n417), .B(KEYINPUT75), .ZN(n479) );
  NAND2_X1 U426 ( .A1(n699), .A2(n416), .ZN(n417) );
  INV_X1 U427 ( .A(G237), .ZN(n416) );
  XNOR2_X1 U428 ( .A(n412), .B(n364), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n411), .B(KEYINPUT98), .ZN(n412) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n411) );
  XNOR2_X1 U431 ( .A(G143), .B(G131), .ZN(n410) );
  XOR2_X1 U432 ( .A(KEYINPUT99), .B(G140), .Z(n415) );
  XNOR2_X1 U433 ( .A(n355), .B(G122), .ZN(n414) );
  XOR2_X1 U434 ( .A(G104), .B(G107), .Z(n454) );
  XOR2_X1 U435 ( .A(G140), .B(KEYINPUT69), .Z(n463) );
  XOR2_X1 U436 ( .A(KEYINPUT104), .B(n532), .Z(n533) );
  NOR2_X1 U437 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U438 ( .A(KEYINPUT5), .B(G113), .Z(n409) );
  XNOR2_X1 U439 ( .A(n451), .B(n450), .ZN(n706) );
  XNOR2_X1 U440 ( .A(n449), .B(G131), .ZN(n450) );
  XOR2_X1 U441 ( .A(G137), .B(KEYINPUT70), .Z(n449) );
  XNOR2_X1 U442 ( .A(G128), .B(G137), .ZN(n464) );
  XNOR2_X1 U443 ( .A(G110), .B(KEYINPUT24), .ZN(n467) );
  XOR2_X1 U444 ( .A(KEYINPUT23), .B(KEYINPUT71), .Z(n468) );
  XNOR2_X1 U445 ( .A(G902), .B(KEYINPUT15), .ZN(n624) );
  XNOR2_X1 U446 ( .A(n362), .B(n452), .ZN(n444) );
  XNOR2_X1 U447 ( .A(n442), .B(n443), .ZN(n362) );
  XNOR2_X1 U448 ( .A(n360), .B(n448), .ZN(n573) );
  XNOR2_X1 U449 ( .A(n406), .B(KEYINPUT73), .ZN(n405) );
  INV_X1 U450 ( .A(KEYINPUT39), .ZN(n406) );
  INV_X1 U451 ( .A(KEYINPUT19), .ZN(n367) );
  XNOR2_X1 U452 ( .A(n571), .B(n348), .ZN(n599) );
  XNOR2_X1 U453 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U454 ( .A(n633), .B(KEYINPUT59), .ZN(n634) );
  NOR2_X1 U455 ( .A1(n610), .A2(n606), .ZN(n598) );
  XNOR2_X1 U456 ( .A(n373), .B(n349), .ZN(n721) );
  INV_X1 U457 ( .A(KEYINPUT32), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n351), .B(n350), .ZN(n535) );
  INV_X1 U459 ( .A(KEYINPUT88), .ZN(n350) );
  NOR2_X1 U460 ( .A1(n533), .A2(KEYINPUT22), .ZN(n344) );
  XOR2_X1 U461 ( .A(n468), .B(n467), .Z(n345) );
  XOR2_X1 U462 ( .A(n415), .B(n414), .Z(n346) );
  AND2_X1 U463 ( .A1(n647), .A2(n536), .ZN(n347) );
  NAND2_X1 U464 ( .A1(n539), .A2(n344), .ZN(n398) );
  XOR2_X1 U465 ( .A(KEYINPUT1), .B(KEYINPUT68), .Z(n348) );
  INV_X1 U466 ( .A(KEYINPUT22), .ZN(n401) );
  XOR2_X1 U467 ( .A(n396), .B(KEYINPUT67), .Z(n349) );
  NAND2_X1 U468 ( .A1(n358), .A2(n398), .ZN(n351) );
  XNOR2_X2 U469 ( .A(n352), .B(KEYINPUT103), .ZN(n659) );
  NAND2_X1 U470 ( .A1(n544), .A2(n502), .ZN(n352) );
  NAND2_X1 U471 ( .A1(n709), .A2(n700), .ZN(n623) );
  NOR2_X2 U472 ( .A1(n381), .A2(n374), .ZN(n709) );
  NAND2_X1 U473 ( .A1(n600), .A2(n359), .ZN(n669) );
  NAND2_X1 U474 ( .A1(n604), .A2(n605), .ZN(n354) );
  XNOR2_X1 U475 ( .A(n548), .B(KEYINPUT44), .ZN(n366) );
  BUF_X1 U476 ( .A(G116), .Z(n356) );
  XNOR2_X1 U477 ( .A(n541), .B(n542), .ZN(n389) );
  NAND2_X1 U478 ( .A1(n366), .A2(n347), .ZN(n365) );
  XNOR2_X1 U479 ( .A(n365), .B(KEYINPUT45), .ZN(n700) );
  BUF_X1 U480 ( .A(n592), .Z(n357) );
  NAND2_X1 U481 ( .A1(n535), .A2(n537), .ZN(n647) );
  XNOR2_X1 U482 ( .A(n425), .B(n426), .ZN(n431) );
  XNOR2_X2 U483 ( .A(n361), .B(n489), .ZN(n540) );
  INV_X1 U484 ( .A(n659), .ZN(n662) );
  NAND2_X1 U485 ( .A1(n659), .A2(n593), .ZN(n594) );
  AND2_X1 U486 ( .A1(n399), .A2(n372), .ZN(n371) );
  NOR2_X2 U487 ( .A1(n400), .A2(n402), .ZN(n399) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n681) );
  INV_X1 U489 ( .A(n434), .ZN(n364) );
  NOR2_X2 U490 ( .A1(n572), .A2(n571), .ZN(n579) );
  NAND2_X1 U491 ( .A1(n379), .A2(n375), .ZN(n374) );
  NAND2_X1 U492 ( .A1(n592), .A2(n596), .ZN(n368) );
  XNOR2_X2 U493 ( .A(n369), .B(n408), .ZN(n592) );
  NAND2_X1 U494 ( .A1(n641), .A2(n624), .ZN(n369) );
  NAND2_X1 U495 ( .A1(n399), .A2(n595), .ZN(n370) );
  NAND2_X1 U496 ( .A1(n371), .A2(n398), .ZN(n373) );
  AND2_X1 U497 ( .A1(n538), .A2(n595), .ZN(n372) );
  NAND2_X1 U498 ( .A1(n398), .A2(n399), .ZN(n546) );
  NAND2_X1 U499 ( .A1(n382), .A2(n380), .ZN(n379) );
  NOR2_X1 U500 ( .A1(n382), .A2(KEYINPUT87), .ZN(n381) );
  NAND2_X1 U501 ( .A1(n561), .A2(n596), .ZN(n503) );
  NOR2_X2 U502 ( .A1(n580), .A2(n524), .ZN(n525) );
  XNOR2_X2 U503 ( .A(n391), .B(n390), .ZN(n571) );
  XNOR2_X2 U504 ( .A(n393), .B(KEYINPUT66), .ZN(n441) );
  XNOR2_X2 U505 ( .A(G143), .B(G128), .ZN(n393) );
  NAND2_X1 U506 ( .A1(n394), .A2(G472), .ZN(n628) );
  NAND2_X1 U507 ( .A1(n394), .A2(G210), .ZN(n643) );
  NAND2_X1 U508 ( .A1(n394), .A2(G475), .ZN(n635) );
  NAND2_X1 U509 ( .A1(n394), .A2(G469), .ZN(n677) );
  NAND2_X1 U510 ( .A1(n394), .A2(G478), .ZN(n682) );
  NAND2_X1 U511 ( .A1(n394), .A2(G217), .ZN(n686) );
  AND2_X2 U512 ( .A1(n627), .A2(n626), .ZN(n394) );
  XNOR2_X2 U513 ( .A(KEYINPUT4), .B(G146), .ZN(n708) );
  INV_X1 U514 ( .A(n721), .ZN(n395) );
  XNOR2_X2 U515 ( .A(n525), .B(KEYINPUT0), .ZN(n539) );
  INV_X1 U516 ( .A(n539), .ZN(n534) );
  NOR2_X1 U517 ( .A1(n539), .A2(n401), .ZN(n400) );
  NAND2_X1 U518 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X2 U519 ( .A(n478), .B(n477), .ZN(n565) );
  XNOR2_X1 U520 ( .A(n403), .B(n345), .ZN(n470) );
  NAND2_X1 U521 ( .A1(n469), .A2(G221), .ZN(n403) );
  XNOR2_X2 U522 ( .A(n407), .B(n405), .ZN(n612) );
  NAND2_X1 U523 ( .A1(n588), .A2(n561), .ZN(n407) );
  XNOR2_X1 U524 ( .A(n677), .B(n676), .ZN(n679) );
  XNOR2_X1 U525 ( .A(n643), .B(n642), .ZN(n644) );
  AND2_X1 U526 ( .A1(G210), .A2(n447), .ZN(n408) );
  INV_X1 U527 ( .A(KEYINPUT65), .ZN(n576) );
  XNOR2_X1 U528 ( .A(n482), .B(n409), .ZN(n483) );
  XNOR2_X1 U529 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U530 ( .A(G472), .ZN(n486) );
  XNOR2_X1 U531 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U532 ( .A(n346), .B(n418), .ZN(n419) );
  XNOR2_X1 U533 ( .A(n458), .B(n459), .ZN(n672) );
  XNOR2_X1 U534 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U537 ( .A(n637), .B(KEYINPUT60), .ZN(n638) );
  XNOR2_X1 U538 ( .A(n619), .B(n618), .ZN(G75) );
  XOR2_X1 U539 ( .A(n410), .B(n462), .Z(n413) );
  XOR2_X1 U540 ( .A(G113), .B(G104), .Z(n434) );
  NAND2_X1 U541 ( .A1(G214), .A2(n479), .ZN(n418) );
  XOR2_X1 U542 ( .A(KEYINPUT101), .B(KEYINPUT13), .Z(n422) );
  XNOR2_X1 U543 ( .A(KEYINPUT100), .B(G475), .ZN(n421) );
  XNOR2_X1 U544 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U545 ( .A(G122), .B(G107), .Z(n433) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(n433), .Z(n426) );
  XNOR2_X1 U547 ( .A(n451), .B(n356), .ZN(n425) );
  XNOR2_X2 U548 ( .A(n699), .B(KEYINPUT64), .ZN(n710) );
  NAND2_X1 U549 ( .A1(n469), .A2(G217), .ZN(n429) );
  XOR2_X1 U550 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n428) );
  NOR2_X1 U551 ( .A1(n681), .A2(G902), .ZN(n432) );
  NAND2_X1 U552 ( .A1(n543), .A2(n544), .ZN(n530) );
  XOR2_X1 U553 ( .A(n434), .B(n433), .Z(n437) );
  XNOR2_X1 U554 ( .A(n482), .B(KEYINPUT16), .ZN(n436) );
  XNOR2_X1 U555 ( .A(n436), .B(n437), .ZN(n690) );
  XNOR2_X1 U556 ( .A(KEYINPUT79), .B(KEYINPUT18), .ZN(n438) );
  XNOR2_X1 U557 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U558 ( .A(n690), .B(n440), .ZN(n445) );
  XNOR2_X1 U559 ( .A(KEYINPUT92), .B(G110), .ZN(n693) );
  NAND2_X1 U560 ( .A1(G224), .A2(n710), .ZN(n443) );
  XNOR2_X1 U561 ( .A(n445), .B(n444), .ZN(n641) );
  XOR2_X1 U562 ( .A(KEYINPUT74), .B(n446), .Z(n447) );
  NAND2_X1 U563 ( .A1(n447), .A2(G214), .ZN(n596) );
  XNOR2_X1 U564 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n448) );
  XOR2_X1 U565 ( .A(KEYINPUT89), .B(KEYINPUT33), .Z(n489) );
  XNOR2_X1 U566 ( .A(n706), .B(n463), .ZN(n459) );
  XOR2_X1 U567 ( .A(n452), .B(n693), .Z(n457) );
  NAND2_X1 U568 ( .A1(G227), .A2(n710), .ZN(n453) );
  XNOR2_X1 U569 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U570 ( .A(n455), .B(KEYINPUT77), .ZN(n456) );
  NAND2_X1 U571 ( .A1(n624), .A2(G234), .ZN(n460) );
  XNOR2_X1 U572 ( .A(n460), .B(KEYINPUT20), .ZN(n472) );
  NAND2_X1 U573 ( .A1(n472), .A2(G221), .ZN(n461) );
  XNOR2_X1 U574 ( .A(KEYINPUT21), .B(n461), .ZN(n531) );
  XNOR2_X1 U575 ( .A(n463), .B(n462), .ZN(n705) );
  XOR2_X1 U576 ( .A(G119), .B(n355), .Z(n465) );
  XNOR2_X1 U577 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U578 ( .A(n705), .B(n466), .ZN(n471) );
  NOR2_X1 U579 ( .A1(n685), .A2(G902), .ZN(n478) );
  AND2_X1 U580 ( .A1(n472), .A2(G217), .ZN(n476) );
  XOR2_X1 U581 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n474) );
  XNOR2_X1 U582 ( .A(KEYINPUT96), .B(KEYINPUT76), .ZN(n473) );
  XNOR2_X1 U583 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U584 ( .A1(G210), .A2(n479), .ZN(n481) );
  XNOR2_X1 U585 ( .A(n480), .B(n481), .ZN(n484) );
  XOR2_X1 U586 ( .A(n706), .B(n485), .Z(n620) );
  NOR2_X1 U587 ( .A1(n620), .A2(G902), .ZN(n487) );
  BUF_X1 U588 ( .A(n555), .Z(n568) );
  XNOR2_X1 U589 ( .A(n555), .B(KEYINPUT6), .ZN(n595) );
  NOR2_X1 U590 ( .A1(n518), .A2(n595), .ZN(n488) );
  NAND2_X1 U591 ( .A1(n573), .A2(n540), .ZN(n515) );
  XNOR2_X1 U592 ( .A(n490), .B(KEYINPUT94), .ZN(n491) );
  XNOR2_X1 U593 ( .A(KEYINPUT14), .B(n491), .ZN(n520) );
  NAND2_X1 U594 ( .A1(G952), .A2(n520), .ZN(n519) );
  INV_X1 U595 ( .A(n519), .ZN(n513) );
  XNOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT52), .ZN(n511) );
  INV_X1 U597 ( .A(n531), .ZN(n564) );
  XNOR2_X1 U598 ( .A(n565), .B(KEYINPUT105), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n564), .A2(n537), .ZN(n492) );
  XNOR2_X1 U600 ( .A(n492), .B(KEYINPUT49), .ZN(n496) );
  INV_X1 U601 ( .A(n599), .ZN(n607) );
  NAND2_X1 U602 ( .A1(n607), .A2(n518), .ZN(n493) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(n493), .Z(n494) );
  NOR2_X1 U604 ( .A1(n568), .A2(n494), .ZN(n495) );
  NAND2_X1 U605 ( .A1(n496), .A2(n495), .ZN(n498) );
  NOR2_X1 U606 ( .A1(n607), .A2(n518), .ZN(n497) );
  NAND2_X1 U607 ( .A1(n568), .A2(n497), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n498), .A2(n527), .ZN(n499) );
  XOR2_X1 U609 ( .A(KEYINPUT51), .B(n499), .Z(n500) );
  NAND2_X1 U610 ( .A1(n573), .A2(n500), .ZN(n509) );
  NOR2_X1 U611 ( .A1(n561), .A2(n596), .ZN(n501) );
  NOR2_X1 U612 ( .A1(n530), .A2(n501), .ZN(n506) );
  INV_X1 U613 ( .A(n543), .ZN(n502) );
  NOR2_X1 U614 ( .A1(n544), .A2(n502), .ZN(n655) );
  NOR2_X1 U615 ( .A1(n586), .A2(n503), .ZN(n504) );
  XOR2_X1 U616 ( .A(KEYINPUT115), .B(n504), .Z(n505) );
  OR2_X1 U617 ( .A1(n506), .A2(n505), .ZN(n507) );
  NAND2_X1 U618 ( .A1(n540), .A2(n507), .ZN(n508) );
  NAND2_X1 U619 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U620 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U621 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U622 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U623 ( .A(n516), .B(KEYINPUT117), .ZN(n517) );
  NAND2_X1 U624 ( .A1(n517), .A2(n699), .ZN(n617) );
  NOR2_X1 U625 ( .A1(n343), .A2(n519), .ZN(n553) );
  NAND2_X1 U626 ( .A1(G902), .A2(n520), .ZN(n549) );
  INV_X1 U627 ( .A(n549), .ZN(n521) );
  NOR2_X1 U628 ( .A1(G898), .A2(n699), .ZN(n695) );
  NAND2_X1 U629 ( .A1(n521), .A2(n695), .ZN(n522) );
  XNOR2_X1 U630 ( .A(KEYINPUT95), .B(n522), .ZN(n523) );
  NOR2_X1 U631 ( .A1(n553), .A2(n523), .ZN(n524) );
  NOR2_X1 U632 ( .A1(n568), .A2(n534), .ZN(n526) );
  NAND2_X1 U633 ( .A1(n559), .A2(n526), .ZN(n649) );
  NOR2_X1 U634 ( .A1(n527), .A2(n534), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n528), .B(KEYINPUT31), .ZN(n665) );
  NAND2_X1 U636 ( .A1(n649), .A2(n665), .ZN(n529) );
  XOR2_X1 U637 ( .A(n586), .B(KEYINPUT84), .Z(n582) );
  NAND2_X1 U638 ( .A1(n529), .A2(n582), .ZN(n536) );
  NOR2_X1 U639 ( .A1(n607), .A2(n537), .ZN(n538) );
  XOR2_X1 U640 ( .A(KEYINPUT34), .B(KEYINPUT80), .Z(n542) );
  NAND2_X1 U641 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U642 ( .A1(n544), .A2(n543), .ZN(n587) );
  OR2_X1 U643 ( .A1(n568), .A2(n359), .ZN(n545) );
  NOR2_X1 U644 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U645 ( .A1(n565), .A2(n547), .ZN(n654) );
  XOR2_X1 U646 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n563) );
  NOR2_X1 U647 ( .A1(n710), .A2(n549), .ZN(n550) );
  XOR2_X1 U648 ( .A(KEYINPUT106), .B(n550), .Z(n551) );
  NOR2_X1 U649 ( .A1(G900), .A2(n551), .ZN(n552) );
  NOR2_X1 U650 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U651 ( .A(KEYINPUT81), .B(n554), .Z(n567) );
  XOR2_X1 U652 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n557) );
  NAND2_X1 U653 ( .A1(n555), .A2(n596), .ZN(n556) );
  XNOR2_X1 U654 ( .A(n557), .B(n556), .ZN(n558) );
  NOR2_X2 U655 ( .A1(n567), .A2(n560), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n659), .A2(n612), .ZN(n562) );
  XNOR2_X1 U657 ( .A(n563), .B(n562), .ZN(n718) );
  XOR2_X1 U658 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n575) );
  NAND2_X1 U659 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U660 ( .A1(n593), .A2(n568), .ZN(n570) );
  XNOR2_X1 U661 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n569) );
  XOR2_X1 U662 ( .A(n570), .B(n569), .Z(n572) );
  NAND2_X1 U663 ( .A1(n579), .A2(n573), .ZN(n574) );
  XNOR2_X1 U664 ( .A(n575), .B(n574), .ZN(n719) );
  XNOR2_X1 U665 ( .A(n578), .B(n577), .ZN(n605) );
  INV_X1 U666 ( .A(n579), .ZN(n581) );
  XOR2_X1 U667 ( .A(n660), .B(KEYINPUT47), .Z(n585) );
  INV_X1 U668 ( .A(n582), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n660), .A2(n583), .ZN(n584) );
  AND2_X1 U670 ( .A1(n585), .A2(n584), .ZN(n603) );
  NAND2_X1 U671 ( .A1(KEYINPUT47), .A2(n586), .ZN(n590) );
  AND2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n357), .A2(n589), .ZN(n658) );
  NAND2_X1 U674 ( .A1(n590), .A2(n658), .ZN(n591) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT83), .ZN(n601) );
  INV_X1 U676 ( .A(n357), .ZN(n610) );
  NOR2_X1 U677 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n597), .A2(n596), .ZN(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT36), .B(n598), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n601), .A2(n669), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U682 ( .A(KEYINPUT107), .B(n606), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(KEYINPUT43), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n671) );
  NAND2_X1 U686 ( .A1(n655), .A2(n612), .ZN(n670) );
  BUF_X2 U687 ( .A(n623), .Z(n621) );
  NOR2_X1 U688 ( .A1(KEYINPUT82), .A2(n621), .ZN(n615) );
  NAND2_X1 U689 ( .A1(KEYINPUT82), .A2(n621), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(KEYINPUT2), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n618) );
  XOR2_X1 U694 ( .A(n620), .B(KEYINPUT62), .Z(n629) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT2), .ZN(n627) );
  INV_X1 U696 ( .A(KEYINPUT86), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(n631) );
  NOR2_X1 U699 ( .A1(G952), .A2(n710), .ZN(n630) );
  XOR2_X1 U700 ( .A(KEYINPUT91), .B(n630), .Z(n689) );
  INV_X1 U701 ( .A(n689), .ZN(n678) );
  NAND2_X1 U702 ( .A1(n631), .A2(n678), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U704 ( .A1(n636), .A2(n678), .ZN(n639) );
  INV_X1 U705 ( .A(KEYINPUT122), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n639), .B(n638), .ZN(G60) );
  XOR2_X1 U707 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n640) );
  NAND2_X1 U708 ( .A1(n644), .A2(n678), .ZN(n646) );
  INV_X1 U709 ( .A(KEYINPUT56), .ZN(n645) );
  XNOR2_X1 U710 ( .A(n646), .B(n645), .ZN(G51) );
  XNOR2_X1 U711 ( .A(G101), .B(n647), .ZN(G3) );
  NOR2_X1 U712 ( .A1(n662), .A2(n649), .ZN(n648) );
  XOR2_X1 U713 ( .A(G104), .B(n648), .Z(G6) );
  INV_X1 U714 ( .A(n655), .ZN(n666) );
  NOR2_X1 U715 ( .A1(n666), .A2(n649), .ZN(n651) );
  XNOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(G107), .B(n652), .ZN(G9) );
  XOR2_X1 U719 ( .A(G110), .B(KEYINPUT113), .Z(n653) );
  XNOR2_X1 U720 ( .A(n654), .B(n653), .ZN(G12) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n657) );
  NAND2_X1 U722 ( .A1(n660), .A2(n655), .ZN(n656) );
  XNOR2_X1 U723 ( .A(n657), .B(n656), .ZN(G30) );
  XNOR2_X1 U724 ( .A(G143), .B(n658), .ZN(G45) );
  NAND2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U726 ( .A(n661), .B(n355), .ZN(G48) );
  NOR2_X1 U727 ( .A1(n662), .A2(n665), .ZN(n663) );
  XOR2_X1 U728 ( .A(G113), .B(n663), .Z(n664) );
  XNOR2_X1 U729 ( .A(KEYINPUT114), .B(n664), .ZN(G15) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U731 ( .A(n356), .B(n667), .Z(G18) );
  XOR2_X1 U732 ( .A(G125), .B(KEYINPUT37), .Z(n668) );
  XNOR2_X1 U733 ( .A(n669), .B(n668), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G134), .B(n670), .ZN(G36) );
  XNOR2_X1 U735 ( .A(G140), .B(n671), .ZN(G42) );
  XOR2_X1 U736 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n674) );
  XNOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n680), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U741 ( .A(KEYINPUT123), .B(n681), .ZN(n683) );
  XOR2_X1 U742 ( .A(n683), .B(n682), .Z(n684) );
  NOR2_X1 U743 ( .A1(n689), .A2(n684), .ZN(G63) );
  XNOR2_X1 U744 ( .A(n685), .B(KEYINPUT124), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(G66) );
  XNOR2_X1 U747 ( .A(n690), .B(G101), .ZN(n691) );
  XNOR2_X1 U748 ( .A(n691), .B(KEYINPUT126), .ZN(n692) );
  XOR2_X1 U749 ( .A(n693), .B(n692), .Z(n694) );
  NOR2_X1 U750 ( .A1(n695), .A2(n694), .ZN(n704) );
  XOR2_X1 U751 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n697) );
  NAND2_X1 U752 ( .A1(G224), .A2(n343), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U754 ( .A1(n698), .A2(G898), .ZN(n702) );
  NAND2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(G69) );
  XOR2_X1 U758 ( .A(n706), .B(n705), .Z(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(n712) );
  XOR2_X1 U760 ( .A(n709), .B(n712), .Z(n711) );
  NAND2_X1 U761 ( .A1(n711), .A2(n710), .ZN(n717) );
  XNOR2_X1 U762 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n713), .A2(G900), .ZN(n714) );
  XOR2_X1 U764 ( .A(KEYINPUT127), .B(n714), .Z(n715) );
  NAND2_X1 U765 ( .A1(n343), .A2(n715), .ZN(n716) );
  NAND2_X1 U766 ( .A1(n717), .A2(n716), .ZN(G72) );
  XOR2_X1 U767 ( .A(n718), .B(G131), .Z(G33) );
  XOR2_X1 U768 ( .A(n719), .B(G137), .Z(G39) );
  XNOR2_X1 U769 ( .A(n720), .B(G122), .ZN(G24) );
  XOR2_X1 U770 ( .A(n721), .B(G119), .Z(G21) );
endmodule

