//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT70), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT70), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(G113gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G120gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(KEYINPUT71), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G113gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n214), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n218), .B1(new_n207), .B2(G134gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n202), .A2(G127gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n220), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G141gat), .B(G148gat), .Z(new_n231));
  INV_X1    g030(.A(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G162gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(KEYINPUT2), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G141gat), .B(G148gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n234), .C1(new_n239), .C2(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT4), .B1(new_n230), .B2(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n212), .A2(new_n219), .B1(new_n225), .B2(new_n228), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n238), .A2(new_n240), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n238), .A2(new_n240), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n230), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n255));
  OR3_X1    g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n244), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n225), .A2(new_n228), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n206), .A2(new_n211), .B1(new_n217), .B2(new_n218), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n241), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n230), .A2(KEYINPUT83), .A3(new_n241), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n254), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n242), .A2(new_n266), .A3(new_n246), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT81), .A4(new_n245), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n268), .A3(new_n253), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT82), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n251), .A2(new_n253), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n242), .A2(new_n246), .A3(new_n266), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n268), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT85), .B(new_n265), .C1(new_n270), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(new_n265), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n256), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT0), .ZN(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G85gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n280), .B2(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(new_n256), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n277), .A2(new_n278), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT85), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n277), .A2(new_n276), .A3(new_n278), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(new_n284), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n286), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n296));
  XOR2_X1   g095(.A(G197gat), .B(G204gat), .Z(new_n297));
  NAND2_X1  g096(.A1(G211gat), .A2(G218gat), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT74), .B(KEYINPUT22), .Z(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(G211gat), .A2(G218gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n298), .B(new_n301), .C1(new_n299), .C2(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT75), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT25), .B1(new_n307), .B2(KEYINPUT23), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT68), .B(G183gat), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n309), .A2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT24), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n308), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT23), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G169gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(KEYINPUT67), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n325), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n317), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331));
  INV_X1    g130(.A(new_n307), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n333), .B2(new_n332), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n313), .A2(new_n315), .B1(new_n311), .B2(new_n312), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  NOR2_X1   g137(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n309), .B2(KEYINPUT27), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n340), .B2(G190gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n324), .B1(KEYINPUT26), .B2(new_n332), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n346), .A3(new_n320), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n345), .A2(new_n347), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n330), .A2(new_n337), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n350), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT77), .B(new_n350), .C1(new_n349), .C2(new_n353), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n306), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OR3_X1    g159(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n350), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n349), .B2(new_n350), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n350), .B1(new_n349), .B2(KEYINPUT29), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n305), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n358), .B2(KEYINPUT78), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n296), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n357), .ZN(new_n372));
  INV_X1    g171(.A(new_n306), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n376), .A2(new_n359), .A3(KEYINPUT80), .A4(new_n365), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n360), .A2(new_n366), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n370), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n376), .A2(new_n359), .A3(new_n365), .A4(new_n370), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n295), .A2(new_n378), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G22gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n250), .A2(new_n352), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n373), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n305), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n249), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n241), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n305), .B1(new_n250), .B2(new_n352), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT3), .B1(new_n305), .B2(new_n352), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n393), .A2(KEYINPUT86), .B1(new_n394), .B2(new_n244), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n393), .A2(KEYINPUT86), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n386), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n385), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(new_n385), .A3(new_n397), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G78gat), .B(G106gat), .Z(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n399), .A2(new_n405), .A3(new_n400), .A4(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT72), .B(G71gat), .ZN(new_n410));
  INV_X1    g209(.A(G99gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G15gat), .B(G43gat), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n330), .A2(new_n337), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n344), .A2(new_n348), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n243), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n349), .A2(new_n230), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n419), .B(KEYINPUT64), .Z(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(KEYINPUT65), .Z(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(KEYINPUT32), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n417), .A2(new_n418), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT34), .B1(new_n429), .B2(new_n420), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(new_n418), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n421), .A2(KEYINPUT34), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n426), .A3(new_n427), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n434), .A2(new_n426), .A3(new_n427), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n427), .B2(new_n426), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n384), .A2(new_n409), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT89), .B1(new_n293), .B2(new_n284), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT6), .B1(new_n293), .B2(new_n284), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n280), .A2(new_n448), .A3(new_n285), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT90), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n286), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n294), .A2(KEYINPUT90), .A3(KEYINPUT6), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .A4(new_n381), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n367), .A2(KEYINPUT37), .A3(new_n377), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n370), .B1(new_n379), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n363), .A2(new_n364), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n460), .A2(new_n305), .B1(new_n372), .B2(new_n373), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT38), .B1(new_n461), .B2(KEYINPUT37), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n454), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n252), .A2(new_n254), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n252), .A2(KEYINPUT88), .A3(new_n254), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n262), .A2(new_n263), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n253), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n284), .B(new_n472), .C1(new_n473), .C2(KEYINPUT39), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT40), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n475), .A2(new_n446), .A3(new_n449), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n409), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n445), .B1(new_n464), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n436), .A2(new_n439), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n409), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n295), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n286), .B(KEYINPUT90), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n450), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n409), .A2(new_n483), .A3(KEYINPUT35), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n482), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G57gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G64gat), .ZN(new_n494));
  INV_X1    g293(.A(G64gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G57gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(G71gat), .A2(G78gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G71gat), .A2(G78gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n497), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(KEYINPUT97), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT97), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(G71gat), .A3(G78gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT96), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(G71gat), .B2(G78gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n510), .A3(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n503), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT98), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G183gat), .B(G211gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n385), .A2(G15gat), .ZN(new_n524));
  INV_X1    g323(.A(G15gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(G1gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT16), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n528), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n525), .A2(G22gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n385), .A2(G15gat), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT93), .B(new_n527), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G8gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n538), .A3(new_n528), .ZN(new_n539));
  AOI21_X1  g338(.A(G1gat), .B1(new_n524), .B2(new_n526), .ZN(new_n540));
  AND2_X1   g339(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n537), .A2(G8gat), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n517), .B2(new_n516), .ZN(new_n544));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n544), .B(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n523), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n523), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G43gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G50gat), .ZN(new_n553));
  INV_X1    g352(.A(G50gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G43gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT15), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G36gat), .ZN(new_n558));
  AND2_X1   g357(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT15), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n552), .A2(KEYINPUT91), .A3(G50gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n552), .B2(G50gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n554), .A2(G43gat), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n565), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n557), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n556), .B1(new_n561), .B2(new_n563), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT17), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n564), .A2(new_n557), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT15), .B1(new_n569), .B2(KEYINPUT91), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n555), .A3(new_n567), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n576), .A2(new_n577), .B1(new_n561), .B2(new_n563), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n574), .B(new_n575), .C1(new_n578), .C2(new_n557), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT8), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n581), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n580), .ZN(new_n590));
  NOR2_X1   g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n590), .A2(new_n591), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n573), .A2(new_n579), .A3(new_n593), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n571), .A2(new_n572), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n593), .A2(new_n599), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n601), .A2(new_n602), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n611), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT101), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n589), .A2(new_n592), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT10), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n516), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n505), .A2(new_n510), .A3(new_n507), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n510), .B1(new_n505), .B2(new_n507), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n515), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n504), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n602), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n597), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n589), .A2(new_n592), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n628), .B1(new_n633), .B2(new_n516), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n623), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n494), .A2(new_n496), .B1(new_n502), .B2(new_n501), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n512), .B2(new_n513), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n631), .B(new_n632), .C1(new_n641), .C2(new_n504), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(new_n638), .A3(new_n628), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n619), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT100), .B1(new_n636), .B2(new_n638), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT10), .B1(new_n642), .B2(new_n628), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n648), .B(new_n637), .C1(new_n649), .C2(new_n623), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n644), .A2(new_n619), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n650), .A4(new_n651), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n646), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n551), .A2(new_n615), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n573), .A2(new_n543), .A3(new_n579), .ZN(new_n658));
  AOI22_X1  g457(.A1(KEYINPUT93), .A2(new_n540), .B1(new_n529), .B2(KEYINPUT92), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n538), .B1(new_n659), .B2(new_n533), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n542), .A2(new_n539), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n601), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT94), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n575), .B1(new_n578), .B2(new_n557), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n543), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n543), .A2(new_n666), .A3(new_n667), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n662), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n663), .B(KEYINPUT13), .Z(new_n672));
  AOI21_X1  g471(.A(KEYINPUT95), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n662), .ZN(new_n674));
  OAI211_X1 g473(.A(KEYINPUT95), .B(new_n672), .C1(new_n674), .C2(new_n668), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n665), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G113gat), .B(G141gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G197gat), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT11), .B(G169gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT12), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n665), .B(new_n682), .C1(new_n673), .C2(new_n676), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n657), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT103), .B1(new_n492), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n691), .B(new_n688), .C1(new_n481), .C2(new_n491), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n295), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n527), .ZN(G1324gat));
  OAI21_X1  g494(.A(new_n477), .B1(new_n690), .B2(new_n692), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT104), .B(new_n477), .C1(new_n690), .C2(new_n692), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(G8gat), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT16), .B(G8gat), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n696), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n698), .B2(new_n699), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n700), .B(new_n703), .C1(new_n704), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g504(.A1(new_n444), .A2(new_n440), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT106), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n444), .A2(new_n708), .A3(new_n440), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n693), .A2(new_n525), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n525), .B1(new_n693), .B2(new_n483), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT105), .B(new_n525), .C1(new_n693), .C2(new_n483), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(G1326gat));
  NOR2_X1   g516(.A1(new_n693), .A2(new_n479), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n718), .B(new_n719), .Z(G1327gat));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n409), .B1(new_n476), .B2(new_n477), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n458), .A2(new_n462), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n487), .A2(new_n723), .A3(new_n450), .A4(new_n381), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n459), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n707), .A2(new_n709), .B1(new_n384), .B2(new_n409), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n725), .A2(new_n726), .B1(new_n486), .B2(new_n490), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n721), .B1(new_n727), .B2(new_n615), .ZN(new_n728));
  INV_X1    g527(.A(new_n295), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n409), .B1(new_n729), .B2(new_n477), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n706), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n454), .A2(new_n459), .A3(new_n463), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n488), .A2(new_n489), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n734), .A2(new_n482), .B1(KEYINPUT35), .B2(new_n485), .ZN(new_n735));
  OAI211_X1 g534(.A(KEYINPUT44), .B(new_n614), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n654), .A2(new_n655), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n645), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n551), .A2(new_n687), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G29gat), .B1(new_n741), .B2(new_n295), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n492), .A2(new_n614), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n562), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n744), .A2(new_n743), .A3(new_n745), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(G1328gat));
  OAI21_X1  g547(.A(G36gat), .B1(new_n741), .B2(new_n482), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n477), .A2(new_n558), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT46), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(G1329gat));
  NOR2_X1   g552(.A1(new_n483), .A2(G43gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT109), .B1(new_n744), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n615), .B1(new_n481), .B2(new_n491), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n757), .A2(new_n758), .A3(new_n740), .A4(new_n754), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT47), .B1(new_n760), .B2(KEYINPUT108), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n728), .A2(new_n736), .A3(new_n710), .A4(new_n740), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n763), .B(new_n760), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1330gat));
  NAND4_X1  g566(.A1(new_n728), .A2(new_n736), .A3(new_n409), .A4(new_n740), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G50gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n757), .A2(new_n554), .A3(new_n409), .A4(new_n740), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n769), .B(new_n772), .C1(new_n770), .C2(KEYINPUT48), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1331gat));
  NAND2_X1  g575(.A1(new_n725), .A2(new_n726), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n491), .ZN(new_n778));
  INV_X1    g577(.A(new_n551), .ZN(new_n779));
  NOR4_X1   g578(.A1(new_n779), .A2(new_n686), .A3(new_n614), .A4(new_n656), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n783), .A3(new_n780), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n729), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n477), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT49), .B(G64gat), .Z(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n788), .B2(new_n790), .ZN(G1333gat));
  NAND3_X1  g590(.A1(new_n782), .A2(new_n710), .A3(new_n784), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G71gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n483), .A2(G71gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n782), .A2(new_n784), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(KEYINPUT50), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n409), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n551), .A2(new_n686), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n656), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n737), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n295), .ZN(new_n807));
  XNOR2_X1  g606(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n778), .A2(new_n614), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n727), .A2(new_n615), .A3(new_n804), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(KEYINPUT112), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n585), .A3(new_n729), .A4(new_n739), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n807), .A2(new_n815), .ZN(G1336gat));
  OR2_X1    g615(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n482), .A2(new_n656), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(G92gat), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n814), .A2(new_n820), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n728), .A2(new_n736), .A3(new_n477), .A4(new_n805), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G92gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n817), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n615), .B1(new_n777), .B2(new_n491), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n813), .B1(new_n825), .B2(new_n803), .ZN(new_n826));
  NOR4_X1   g625(.A1(new_n727), .A2(new_n615), .A3(new_n804), .A4(new_n808), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n820), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n823), .A2(new_n828), .A3(new_n829), .A4(new_n817), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n824), .A2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n806), .B2(new_n711), .ZN(new_n832));
  INV_X1    g631(.A(new_n483), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n814), .A2(new_n411), .A3(new_n833), .A4(new_n739), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1338gat));
  NOR3_X1   g634(.A1(new_n479), .A2(G106gat), .A3(new_n656), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n728), .A2(new_n736), .A3(new_n409), .A4(new_n805), .ZN(new_n838));
  XOR2_X1   g637(.A(KEYINPUT114), .B(G106gat), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1339gat));
  NAND3_X1  g644(.A1(new_n686), .A2(new_n221), .A3(new_n223), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n636), .B2(new_n638), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n647), .A2(new_n850), .A3(new_n650), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n849), .B(new_n637), .C1(new_n649), .C2(new_n623), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(KEYINPUT115), .A3(new_n619), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT115), .B1(new_n852), .B2(new_n619), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n851), .B(KEYINPUT55), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n738), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n619), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n853), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT55), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT116), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n738), .A4(new_n856), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n863), .A2(new_n686), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n674), .A2(new_n672), .A3(new_n668), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n663), .B1(new_n658), .B2(new_n662), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n870), .B(new_n681), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n681), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT117), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n685), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n739), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n685), .A2(new_n873), .A3(new_n875), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT118), .B1(new_n879), .B2(new_n656), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n615), .B1(new_n869), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n615), .A2(new_n879), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n863), .A3(new_n868), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n551), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n657), .A2(new_n686), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n848), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n877), .B1(new_n876), .B2(new_n739), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n879), .A2(new_n656), .A3(KEYINPUT118), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n863), .A2(new_n686), .A3(new_n868), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n614), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n884), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n779), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n886), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(KEYINPUT119), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n887), .A2(new_n729), .A3(new_n484), .A4(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n482), .B(new_n847), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n894), .A2(KEYINPUT119), .A3(new_n895), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT119), .B1(new_n894), .B2(new_n895), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n902), .A2(new_n903), .A3(new_n409), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n482), .A2(new_n729), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n904), .A2(new_n833), .A3(new_n686), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G113gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1340gat));
  OAI21_X1  g712(.A(new_n482), .B1(new_n899), .B2(new_n900), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(new_n656), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n904), .A2(new_n906), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n483), .A2(new_n213), .A3(new_n656), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n915), .A2(new_n213), .B1(new_n917), .B2(new_n918), .ZN(G1341gat));
  AND2_X1   g718(.A1(new_n208), .A2(new_n210), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n551), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n916), .A2(new_n483), .A3(new_n779), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n914), .A2(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1342gat));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n904), .A2(new_n833), .A3(new_n614), .A4(new_n906), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G134gat), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n482), .A2(new_n203), .A3(new_n205), .A4(new_n614), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n902), .A2(new_n903), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n928), .A2(KEYINPUT120), .A3(new_n729), .A4(new_n484), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n897), .A2(new_n898), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g732(.A(KEYINPUT56), .B(new_n927), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n924), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n927), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(new_n899), .B2(new_n900), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT56), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n931), .A2(new_n932), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n938), .A2(KEYINPUT122), .A3(new_n939), .A4(new_n926), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n935), .A2(new_n940), .ZN(G1343gat));
  INV_X1    g740(.A(G141gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n887), .A2(new_n896), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(new_n295), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n710), .A2(new_n479), .A3(new_n477), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n946), .B2(new_n687), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT57), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n948), .A3(new_n409), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n711), .A2(new_n906), .ZN(new_n950));
  INV_X1    g749(.A(new_n864), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n865), .B1(new_n951), .B2(KEYINPUT123), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(KEYINPUT123), .B2(new_n951), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n686), .A2(new_n738), .A3(new_n856), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n953), .A2(new_n954), .B1(new_n656), .B2(new_n879), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n615), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n551), .B1(new_n956), .B2(new_n884), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n409), .B1(new_n957), .B2(new_n886), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n950), .B1(KEYINPUT57), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n686), .A2(G141gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n947), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT58), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n947), .B(KEYINPUT58), .C1(new_n960), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1344gat));
  INV_X1    g765(.A(new_n946), .ZN(new_n967));
  INV_X1    g766(.A(G148gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(new_n739), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n960), .A2(new_n656), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n970), .A2(KEYINPUT59), .A3(new_n968), .ZN(new_n971));
  XOR2_X1   g770(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n972));
  OAI21_X1  g771(.A(KEYINPUT57), .B1(new_n943), .B2(new_n479), .ZN(new_n973));
  INV_X1    g772(.A(new_n950), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n886), .B(KEYINPUT125), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n883), .A2(new_n738), .A3(new_n856), .A4(new_n866), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n551), .B1(new_n956), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n948), .B(new_n409), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n973), .A2(new_n739), .A3(new_n974), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n972), .B1(new_n979), .B2(G148gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n969), .B1(new_n971), .B2(new_n980), .ZN(G1345gat));
  NAND3_X1  g780(.A1(new_n967), .A2(new_n232), .A3(new_n551), .ZN(new_n982));
  OAI21_X1  g781(.A(G155gat), .B1(new_n960), .B2(new_n779), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1346gat));
  AOI21_X1  g783(.A(G162gat), .B1(new_n967), .B2(new_n614), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n960), .A2(new_n233), .A3(new_n615), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1347gat));
  NAND2_X1  g786(.A1(new_n477), .A2(new_n295), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n988), .A2(new_n483), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n904), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n990), .A2(new_n322), .A3(new_n687), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n943), .A2(new_n729), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n992), .A2(new_n477), .A3(new_n484), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n993), .A2(new_n687), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n991), .B1(new_n994), .B2(new_n322), .ZN(G1348gat));
  OAI21_X1  g794(.A(new_n323), .B1(new_n993), .B2(new_n656), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n739), .A2(G176gat), .ZN(new_n998));
  OR3_X1    g797(.A1(new_n990), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n997), .B1(new_n990), .B2(new_n998), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(G1349gat));
  OAI21_X1  g800(.A(new_n309), .B1(new_n990), .B2(new_n779), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n551), .A2(new_n342), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n993), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g803(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1004), .B(new_n1005), .ZN(G1350gat));
  NAND3_X1  g805(.A1(new_n904), .A2(new_n614), .A3(new_n989), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1007), .A2(new_n1008), .A3(G190gat), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1008), .B1(new_n1007), .B2(G190gat), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n614), .A2(new_n312), .ZN(new_n1012));
  OAI22_X1  g811(.A1(new_n1010), .A2(new_n1011), .B1(new_n993), .B2(new_n1012), .ZN(G1351gat));
  AND2_X1   g812(.A1(new_n973), .A2(new_n978), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n710), .A2(new_n988), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g816(.A(G197gat), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n687), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n710), .A2(new_n479), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n992), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1022), .A2(new_n477), .A3(new_n686), .ZN(new_n1023));
  AOI22_X1  g822(.A1(new_n1017), .A2(new_n1019), .B1(new_n1023), .B2(new_n1018), .ZN(G1352gat));
  NOR2_X1   g823(.A1(new_n819), .A2(G204gat), .ZN(new_n1025));
  AND3_X1   g824(.A1(new_n992), .A2(new_n1020), .A3(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g825(.A(new_n1026), .B(KEYINPUT62), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1014), .A2(new_n739), .A3(new_n1016), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1028), .A2(G204gat), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(new_n1029), .ZN(G1353gat));
  NAND4_X1  g829(.A1(new_n973), .A2(new_n551), .A3(new_n978), .A4(new_n1016), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1031), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(KEYINPUT63), .B1(new_n1031), .B2(G211gat), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1022), .A2(new_n477), .ZN(new_n1034));
  OR2_X1    g833(.A1(new_n779), .A2(G211gat), .ZN(new_n1035));
  OAI22_X1  g834(.A1(new_n1032), .A2(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(G1354gat));
  NAND3_X1  g835(.A1(new_n1014), .A2(new_n614), .A3(new_n1016), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1037), .A2(G218gat), .ZN(new_n1038));
  OR2_X1    g837(.A1(new_n615), .A2(G218gat), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1038), .B1(new_n1034), .B2(new_n1039), .ZN(G1355gat));
endmodule


