//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G137), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n458), .A2(new_n460), .B1(new_n461), .B2(G101), .ZN(new_n462));
  AND2_X1   g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n458), .B2(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n464), .B2(new_n459), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G160));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n458), .A2(KEYINPUT64), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n459), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n459), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n459), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n475), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT65), .Z(G162));
  AND2_X1   g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n458), .A2(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n490), .B(new_n491), .C1(new_n468), .C2(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n458), .B2(new_n490), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(KEYINPUT66), .B(new_n488), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XOR2_X1   g079(.A(new_n504), .B(KEYINPUT68), .Z(new_n505));
  OAI21_X1  g080(.A(G651), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n501), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n507), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT67), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n514), .A2(KEYINPUT67), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n506), .B1(new_n516), .B2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT69), .B(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n501), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n510), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n529), .A2(new_n511), .B1(new_n512), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n533), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n537), .B1(new_n538), .B2(new_n511), .C1(new_n539), .C2(new_n512), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  INV_X1    g121(.A(new_n512), .ZN(new_n547));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n524), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(G91), .A2(new_n547), .B1(new_n550), .B2(G651), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n511), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n508), .A2(new_n509), .ZN(new_n554));
  INV_X1    g129(.A(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(new_n557), .A3(G53), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n551), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  XOR2_X1   g136(.A(G168), .B(KEYINPUT70), .Z(G286));
  OAI21_X1  g137(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n563));
  INV_X1    g138(.A(G87), .ZN(new_n564));
  INV_X1    g139(.A(G49), .ZN(new_n565));
  OAI221_X1 g140(.A(new_n563), .B1(new_n512), .B2(new_n564), .C1(new_n565), .C2(new_n511), .ZN(G288));
  AOI22_X1  g141(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n533), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n547), .A2(G86), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n556), .A2(G48), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  AOI22_X1  g146(.A1(new_n547), .A2(G85), .B1(new_n556), .B2(G47), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n533), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G290));
  INV_X1    g150(.A(G868), .ZN(new_n576));
  NOR2_X1   g151(.A1(G171), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT71), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n547), .A2(G92), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT10), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(KEYINPUT10), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n556), .A2(G54), .ZN(new_n583));
  XOR2_X1   g158(.A(KEYINPUT72), .B(G66), .Z(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(new_n501), .B1(G79), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n585), .B2(new_n533), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n583), .B(KEYINPUT73), .C1(new_n585), .C2(new_n533), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n578), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n578), .B1(new_n592), .B2(G868), .ZN(G321));
  MUX2_X1   g169(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g170(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n592), .B1(new_n597), .B2(G860), .ZN(G148));
  NOR2_X1   g173(.A1(new_n541), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n592), .A2(new_n597), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT74), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n599), .B1(new_n601), .B2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT75), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n474), .A2(G123), .ZN(new_n605));
  OR2_X1    g180(.A1(G99), .A2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n606), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G135), .B2(new_n477), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2096), .ZN(new_n610));
  NAND2_X1  g185(.A1(KEYINPUT76), .A2(G2100), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n458), .A2(new_n461), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  NOR2_X1   g189(.A1(KEYINPUT76), .A2(G2100), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n610), .B(new_n616), .C1(new_n614), .C2(new_n611), .ZN(G156));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(KEYINPUT14), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n626), .B(new_n627), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT78), .Z(new_n632));
  OAI21_X1  g207(.A(G14), .B1(new_n629), .B2(new_n630), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(G401));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2096), .B(G2100), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT79), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n635), .A2(new_n636), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n643), .B(new_n647), .Z(G227));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT81), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n652), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1981), .B(G1986), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT83), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT82), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n665), .B(new_n668), .Z(G229));
  NAND2_X1  g244(.A1(new_n474), .A2(G129), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT94), .ZN(new_n671));
  NAND3_X1  g246(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT26), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n461), .A2(G105), .ZN(new_n674));
  INV_X1    g249(.A(G141), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n673), .B(new_n674), .C1(new_n476), .C2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G29), .ZN(new_n678));
  NOR2_X1   g253(.A1(G29), .A2(G32), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(KEYINPUT95), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(KEYINPUT95), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT27), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT96), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT25), .Z(new_n688));
  INV_X1    g263(.A(G139), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n476), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n693));
  OAI22_X1  g268(.A1(new_n691), .A2(new_n692), .B1(new_n459), .B2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G33), .B(new_n694), .S(G29), .Z(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G2072), .ZN(new_n696));
  NOR2_X1   g271(.A1(G4), .A2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT86), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n591), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1348), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n685), .A2(new_n686), .A3(new_n696), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G26), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n477), .A2(G140), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT89), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(G116), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G2105), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n474), .B2(G128), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n706), .B1(new_n713), .B2(G29), .ZN(new_n714));
  INV_X1    g289(.A(G2067), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G2072), .B2(new_n695), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n699), .A2(G20), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT23), .ZN(new_n719));
  INV_X1    g294(.A(G299), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n699), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT98), .B(G1956), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n699), .A2(G5), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G171), .B2(new_n699), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1961), .ZN(new_n727));
  INV_X1    g302(.A(new_n721), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  INV_X1    g304(.A(G2084), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n731));
  INV_X1    g306(.A(G34), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n733), .A2(new_n704), .A3(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT93), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n736), .B(new_n737), .C1(new_n704), .C2(new_n465), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n609), .A2(G29), .B1(new_n730), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT31), .B(G11), .Z(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n699), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n739), .B(new_n744), .C1(G1966), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n699), .A2(G19), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT87), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n540), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT88), .B(G1341), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n704), .A2(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n704), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2078), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n746), .A2(G1966), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n738), .B2(new_n730), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n747), .A2(new_n752), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n717), .A2(new_n724), .A3(new_n729), .A4(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n704), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n704), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT29), .Z(new_n763));
  AOI211_X1 g338(.A(new_n702), .B(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n760), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  MUX2_X1   g341(.A(G6), .B(G305), .S(G16), .Z(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT85), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  NAND2_X1  g344(.A1(G166), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G22), .ZN(new_n771));
  INV_X1    g346(.A(G1971), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n768), .A2(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n699), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(G288), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n699), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT33), .B(G1976), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n768), .B2(new_n769), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n774), .A2(KEYINPUT34), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT34), .B1(new_n774), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n474), .A2(G119), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n477), .A2(G131), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT84), .B1(G95), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(KEYINPUT84), .A2(G95), .A3(G2105), .ZN(new_n787));
  OAI221_X1 g362(.A(G2104), .B1(G107), .B2(new_n459), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n783), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G29), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G25), .B2(G29), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n699), .A2(G24), .ZN(new_n796));
  INV_X1    g371(.A(G290), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n699), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1986), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n794), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n781), .A2(new_n782), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n764), .B(new_n766), .C1(new_n802), .C2(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  XNOR2_X1  g380(.A(KEYINPUT100), .B(G860), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n591), .A2(new_n597), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G55), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n813), .A2(new_n511), .B1(new_n512), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n533), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n540), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n820), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n810), .A2(new_n811), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  AOI211_X1 g402(.A(KEYINPUT101), .B(new_n827), .C1(new_n821), .C2(new_n823), .ZN(new_n828));
  OAI221_X1 g403(.A(new_n806), .B1(KEYINPUT39), .B2(new_n824), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n818), .A2(new_n806), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(G162), .A2(new_n609), .ZN(new_n835));
  NAND2_X1  g410(.A1(G162), .A2(new_n609), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n465), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n465), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n833), .A3(new_n837), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n713), .B(new_n495), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n790), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n677), .B(new_n694), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n474), .A2(G130), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n477), .A2(G142), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n459), .A2(KEYINPUT104), .A3(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT104), .B1(new_n459), .B2(G118), .ZN(new_n850));
  OR2_X1    g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(G2104), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n613), .Z(new_n854));
  AND2_X1   g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n846), .A2(new_n854), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n845), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n845), .B1(new_n856), .B2(new_n855), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n843), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n842), .B(new_n840), .C1(new_n861), .C2(new_n857), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(new_n601), .B(new_n820), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n591), .A2(G299), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n591), .A2(G299), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .A3(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n776), .B(G290), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT105), .ZN(new_n879));
  XNOR2_X1  g454(.A(G303), .B(G305), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(KEYINPUT105), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT42), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n876), .A2(new_n877), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n876), .B2(new_n877), .ZN(new_n887));
  OAI21_X1  g462(.A(G868), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(G868), .B2(new_n818), .ZN(G295));
  OAI21_X1  g464(.A(new_n888), .B1(G868), .B2(new_n818), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n891));
  NOR2_X1   g466(.A1(G171), .A2(G168), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(G286), .B2(G301), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n822), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n820), .B(new_n893), .C1(G301), .C2(G286), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n868), .A3(new_n872), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n874), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n884), .ZN(new_n900));
  INV_X1    g475(.A(new_n884), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(new_n898), .C1(new_n874), .C2(new_n897), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n902), .A3(new_n863), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n863), .A4(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n891), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI211_X1 g485(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(new_n903), .B2(KEYINPUT43), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n910), .A2(new_n911), .B1(new_n913), .B2(new_n916), .ZN(G397));
  OAI21_X1  g492(.A(new_n490), .B1(new_n467), .B2(new_n468), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT4), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n492), .ZN(new_n920));
  AOI21_X1  g495(.A(G1384), .B1(new_n920), .B2(new_n488), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  INV_X1    g500(.A(G40), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n465), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G125), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n469), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G2105), .B1(new_n929), .B2(new_n463), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(KEYINPUT109), .A3(G40), .A4(new_n462), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n677), .B(G1996), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n713), .B(new_n715), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n790), .A2(new_n793), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n790), .A2(new_n793), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1986), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n797), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT110), .Z(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n939), .B2(new_n797), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n933), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT54), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n497), .B2(new_n498), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT111), .B1(new_n946), .B2(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  INV_X1    g523(.A(new_n498), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT66), .B1(new_n920), .B2(new_n488), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n923), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n921), .A2(KEYINPUT45), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n954), .A2(new_n927), .A3(new_n931), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n947), .A2(new_n953), .A3(new_n958), .A4(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G2078), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT125), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G2078), .B1(new_n957), .B2(new_n959), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT125), .B1(new_n966), .B2(KEYINPUT53), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n499), .B2(new_n948), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n921), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n927), .A3(new_n931), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1961), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n927), .A2(new_n931), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(KEYINPUT116), .A3(new_n924), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT116), .B1(new_n975), .B2(new_n924), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n964), .A2(G2078), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G301), .B1(new_n968), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n465), .A2(new_n926), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n924), .A2(new_n954), .A3(new_n984), .A4(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n973), .B2(G1961), .ZN(new_n986));
  AOI211_X1 g561(.A(G171), .B(new_n986), .C1(new_n965), .C2(new_n967), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n945), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n947), .A2(new_n953), .A3(new_n989), .A4(new_n955), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n975), .A2(new_n921), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT58), .B(G1341), .Z(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n990), .A2(KEYINPUT119), .A3(new_n993), .ZN(new_n998));
  AND4_X1   g573(.A1(new_n541), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n540), .B1(new_n994), .B2(new_n995), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n998), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT122), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT56), .B(G2072), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n947), .A2(new_n953), .A3(new_n955), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1956), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n951), .A2(KEYINPUT50), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n927), .B(new_n931), .C1(new_n921), .C2(new_n969), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT57), .B1(new_n559), .B2(KEYINPUT117), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(G299), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1006), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(KEYINPUT61), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(KEYINPUT121), .A3(new_n1016), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1013), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT61), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1004), .A2(new_n1017), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT123), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n592), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1348), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n970), .B2(new_n972), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n932), .A2(new_n922), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n715), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1027), .A2(KEYINPUT118), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT118), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1025), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n592), .A2(new_n1024), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g609(.A(new_n1025), .B1(new_n1024), .B2(new_n592), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT60), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1017), .A2(new_n1004), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1003), .A2(new_n1022), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1030), .A2(new_n1031), .A3(new_n591), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1019), .B1(new_n1040), .B2(new_n1016), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1966), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n978), .B2(new_n979), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n973), .A2(new_n730), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(G168), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(KEYINPUT124), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n527), .B2(new_n523), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1053), .A3(new_n1048), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n957), .A2(new_n772), .A3(new_n959), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(G2090), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  NOR3_X1   g635(.A1(G166), .A2(new_n1060), .A3(new_n1047), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1060), .B1(G166), .B2(new_n1047), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n776), .A2(G1976), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n991), .A2(G8), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1028), .A2(new_n1047), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1068), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G305), .A2(G1981), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n568), .A2(new_n569), .A3(new_n1076), .A4(new_n570), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1074), .A2(KEYINPUT52), .B1(new_n1080), .B2(new_n1073), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1072), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n973), .A2(new_n760), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1047), .B1(new_n1056), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1055), .A2(new_n1067), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n963), .B1(new_n962), .B2(new_n964), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n966), .A2(KEYINPUT125), .A3(KEYINPUT53), .ZN(new_n1089));
  OAI211_X1 g664(.A(G301), .B(new_n982), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n986), .B1(new_n965), .B2(new_n967), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(KEYINPUT54), .C1(G301), .C2(new_n1091), .ZN(new_n1092));
  AND4_X1   g667(.A1(new_n988), .A2(new_n1042), .A3(new_n1087), .A4(new_n1092), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1047), .B(G286), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1067), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT63), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1094), .A2(KEYINPUT63), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1086), .B(new_n1098), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1067), .A2(new_n1086), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1050), .A2(new_n1103), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1101), .A2(new_n983), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1073), .B(KEYINPUT115), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1080), .A2(new_n1073), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(new_n1069), .A3(new_n776), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(new_n1077), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1082), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1100), .A2(new_n1105), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n944), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n935), .A2(new_n677), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT46), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n933), .A2(new_n989), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n933), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1116), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT126), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT47), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1121), .B(KEYINPUT127), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT47), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n934), .A2(new_n935), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1128), .A2(new_n936), .B1(G2067), .B2(new_n713), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n938), .A2(new_n933), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n941), .A2(new_n933), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT48), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n933), .A2(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1125), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1114), .A2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g710(.A(G319), .ZN(new_n1137));
  NOR2_X1   g711(.A1(G227), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g712(.A(new_n1138), .B1(new_n632), .B2(new_n633), .ZN(new_n1139));
  NOR2_X1   g713(.A1(G229), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n1140), .A2(new_n864), .A3(new_n908), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


