

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(n716), .B(n715), .ZN(n723) );
  XOR2_X1 U553 ( .A(KEYINPUT27), .B(n705), .Z(n519) );
  INV_X1 U554 ( .A(KEYINPUT99), .ZN(n707) );
  XNOR2_X1 U555 ( .A(KEYINPUT29), .B(KEYINPUT100), .ZN(n715) );
  NOR2_X1 U556 ( .A1(n731), .A2(n730), .ZN(n732) );
  INV_X1 U557 ( .A(n975), .ZN(n758) );
  NAND2_X2 U558 ( .A1(n767), .A2(n693), .ZN(n737) );
  AND2_X1 U559 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X2 U560 ( .A1(G2105), .A2(n540), .ZN(n890) );
  NOR2_X1 U561 ( .A1(G651), .A2(n632), .ZN(n660) );
  NOR2_X1 U562 ( .A1(n545), .A2(n544), .ZN(G164) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NAND2_X1 U564 ( .A1(n660), .A2(G51), .ZN(n520) );
  XNOR2_X1 U565 ( .A(n520), .B(KEYINPUT78), .ZN(n523) );
  INV_X1 U566 ( .A(G651), .ZN(n527) );
  NOR2_X1 U567 ( .A1(G543), .A2(n527), .ZN(n521) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n521), .Z(n654) );
  NAND2_X1 U569 ( .A1(G63), .A2(n654), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U571 ( .A(KEYINPUT6), .B(n524), .ZN(n533) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n656) );
  NAND2_X1 U573 ( .A1(G89), .A2(n656), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n525), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n526), .B(KEYINPUT76), .ZN(n529) );
  NOR2_X1 U576 ( .A1(n632), .A2(n527), .ZN(n652) );
  NAND2_X1 U577 ( .A1(G76), .A2(n652), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U579 ( .A(KEYINPUT5), .B(n530), .ZN(n531) );
  XNOR2_X1 U580 ( .A(KEYINPUT77), .B(n531), .ZN(n532) );
  NOR2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT7), .B(n534), .Z(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U584 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n536) );
  NOR2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XNOR2_X2 U586 ( .A(n536), .B(n535), .ZN(n859) );
  NAND2_X1 U587 ( .A1(n859), .A2(G138), .ZN(n539) );
  INV_X1 U588 ( .A(G2104), .ZN(n540) );
  NAND2_X1 U589 ( .A1(G102), .A2(n890), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT89), .B(n537), .Z(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n545) );
  AND2_X1 U592 ( .A1(n540), .A2(G2105), .ZN(n886) );
  NAND2_X1 U593 ( .A1(n886), .A2(G126), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n541) );
  XOR2_X1 U595 ( .A(KEYINPUT64), .B(n541), .Z(n575) );
  NAND2_X1 U596 ( .A1(G114), .A2(n575), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U598 ( .A(G2451), .B(G2446), .ZN(n555) );
  XOR2_X1 U599 ( .A(G2430), .B(KEYINPUT107), .Z(n547) );
  XNOR2_X1 U600 ( .A(G2454), .B(G2435), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n547), .B(n546), .ZN(n551) );
  XOR2_X1 U602 ( .A(G2438), .B(KEYINPUT106), .Z(n549) );
  XNOR2_X1 U603 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U605 ( .A(n551), .B(n550), .Z(n553) );
  XNOR2_X1 U606 ( .A(G2443), .B(G2427), .ZN(n552) );
  XNOR2_X1 U607 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U608 ( .A(n555), .B(n554), .ZN(n556) );
  AND2_X1 U609 ( .A1(n556), .A2(G14), .ZN(G401) );
  NAND2_X1 U610 ( .A1(G90), .A2(n656), .ZN(n558) );
  NAND2_X1 U611 ( .A1(G77), .A2(n652), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n559), .B(KEYINPUT9), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G64), .A2(n654), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U616 ( .A1(n660), .A2(G52), .ZN(n562) );
  XOR2_X1 U617 ( .A(KEYINPUT68), .B(n562), .Z(n563) );
  NOR2_X1 U618 ( .A1(n564), .A2(n563), .ZN(G171) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U620 ( .A1(n886), .A2(G123), .ZN(n566) );
  XNOR2_X1 U621 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n566), .B(n565), .ZN(n573) );
  NAND2_X1 U623 ( .A1(G99), .A2(n890), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G135), .A2(n859), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n571) );
  BUF_X1 U626 ( .A(n575), .Z(n887) );
  NAND2_X1 U627 ( .A1(G111), .A2(n887), .ZN(n569) );
  XNOR2_X1 U628 ( .A(KEYINPUT81), .B(n569), .ZN(n570) );
  NOR2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n920) );
  XNOR2_X1 U631 ( .A(G2096), .B(n920), .ZN(n574) );
  OR2_X1 U632 ( .A1(G2100), .A2(n574), .ZN(G156) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  INV_X1 U635 ( .A(G57), .ZN(G237) );
  NAND2_X1 U636 ( .A1(G137), .A2(n859), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G113), .A2(n575), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U639 ( .A(KEYINPUT66), .B(n578), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n886), .A2(G125), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G101), .A2(n890), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT23), .B(n579), .Z(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U644 ( .A1(n583), .A2(n582), .ZN(G160) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U646 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U647 ( .A(G223), .B(KEYINPUT71), .ZN(n831) );
  NAND2_X1 U648 ( .A1(n831), .A2(G567), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U650 ( .A1(n654), .A2(G56), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT14), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G43), .A2(n660), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n595) );
  NAND2_X1 U654 ( .A1(n656), .A2(G81), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n589), .B(KEYINPUT12), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G68), .A2(n652), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U658 ( .A(KEYINPUT13), .B(n592), .Z(n593) );
  XNOR2_X1 U659 ( .A(KEYINPUT72), .B(n593), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n596), .ZN(n985) );
  INV_X1 U662 ( .A(n985), .ZN(n620) );
  NAND2_X1 U663 ( .A1(n620), .A2(G860), .ZN(G153) );
  XOR2_X1 U664 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT75), .B(n597), .Z(n606) );
  NAND2_X1 U667 ( .A1(G92), .A2(n656), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G79), .A2(n652), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G66), .A2(n654), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G54), .A2(n660), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(KEYINPUT15), .ZN(n966) );
  INV_X1 U675 ( .A(G868), .ZN(n674) );
  NAND2_X1 U676 ( .A1(n966), .A2(n674), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G91), .A2(n656), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G78), .A2(n652), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G65), .A2(n654), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G53), .A2(n660), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT69), .ZN(n976) );
  XNOR2_X1 U686 ( .A(KEYINPUT70), .B(n976), .ZN(G299) );
  NOR2_X1 U687 ( .A1(G299), .A2(G868), .ZN(n615) );
  NOR2_X1 U688 ( .A1(G286), .A2(n674), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(G297) );
  INV_X1 U690 ( .A(G860), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n616), .A2(G559), .ZN(n617) );
  INV_X1 U692 ( .A(n966), .ZN(n902) );
  NAND2_X1 U693 ( .A1(n617), .A2(n902), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(G559), .A2(n966), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n674), .A2(n619), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n620), .A2(G868), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(KEYINPUT79), .B(n623), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G559), .A2(n902), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(n985), .ZN(n672) );
  NOR2_X1 U702 ( .A1(n672), .A2(G860), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G67), .A2(n654), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G55), .A2(n660), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G93), .A2(n656), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G80), .A2(n652), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n675) );
  XOR2_X1 U710 ( .A(n631), .B(n675), .Z(G145) );
  NAND2_X1 U711 ( .A1(G87), .A2(n632), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n633), .B(KEYINPUT82), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G49), .A2(n660), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n654), .A2(n636), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G85), .A2(n656), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G72), .A2(n652), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U721 ( .A(KEYINPUT67), .B(n641), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G60), .A2(n654), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G47), .A2(n660), .ZN(n642) );
  AND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G88), .A2(n656), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G75), .A2(n652), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G62), .A2(n654), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G50), .A2(n660), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U732 ( .A1(n651), .A2(n650), .ZN(G166) );
  NAND2_X1 U733 ( .A1(G73), .A2(n652), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n654), .A2(G61), .ZN(n655) );
  XOR2_X1 U736 ( .A(KEYINPUT83), .B(n655), .Z(n658) );
  NAND2_X1 U737 ( .A1(n656), .A2(G86), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U739 ( .A(KEYINPUT84), .B(n659), .ZN(n663) );
  NAND2_X1 U740 ( .A1(G48), .A2(n660), .ZN(n661) );
  XNOR2_X1 U741 ( .A(KEYINPUT85), .B(n661), .ZN(n662) );
  NOR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(G305) );
  XOR2_X1 U744 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n666) );
  XNOR2_X1 U745 ( .A(G288), .B(n666), .ZN(n667) );
  XOR2_X1 U746 ( .A(n675), .B(n667), .Z(n669) );
  XNOR2_X1 U747 ( .A(G290), .B(G166), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U749 ( .A(G299), .B(n670), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n671), .B(G305), .ZN(n900) );
  XNOR2_X1 U751 ( .A(n672), .B(n900), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n673), .A2(G868), .ZN(n677) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XNOR2_X1 U756 ( .A(n678), .B(KEYINPUT87), .ZN(n679) );
  XNOR2_X1 U757 ( .A(n679), .B(KEYINPUT20), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n680), .A2(G2090), .ZN(n681) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U760 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U762 ( .A1(G120), .A2(G69), .ZN(n683) );
  NOR2_X1 U763 ( .A1(G237), .A2(n683), .ZN(n684) );
  XNOR2_X1 U764 ( .A(KEYINPUT88), .B(n684), .ZN(n685) );
  NAND2_X1 U765 ( .A1(n685), .A2(G108), .ZN(n837) );
  NAND2_X1 U766 ( .A1(n837), .A2(G567), .ZN(n690) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U769 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U770 ( .A1(G96), .A2(n688), .ZN(n836) );
  NAND2_X1 U771 ( .A1(n836), .A2(G2106), .ZN(n689) );
  NAND2_X1 U772 ( .A1(n690), .A2(n689), .ZN(n914) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n691) );
  NOR2_X1 U774 ( .A1(n914), .A2(n691), .ZN(n835) );
  NAND2_X1 U775 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  INV_X1 U777 ( .A(KEYINPUT101), .ZN(n736) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n766) );
  INV_X1 U780 ( .A(n766), .ZN(n693) );
  NAND2_X1 U781 ( .A1(G1348), .A2(n737), .ZN(n695) );
  INV_X1 U782 ( .A(n737), .ZN(n718) );
  NAND2_X1 U783 ( .A1(G2067), .A2(n718), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n702) );
  NOR2_X1 U785 ( .A1(n966), .A2(n702), .ZN(n701) );
  INV_X1 U786 ( .A(G1996), .ZN(n943) );
  NOR2_X1 U787 ( .A1(n737), .A2(n943), .ZN(n696) );
  XOR2_X1 U788 ( .A(n696), .B(KEYINPUT26), .Z(n698) );
  NAND2_X1 U789 ( .A1(n737), .A2(G1341), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n699), .A2(n985), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n704) );
  AND2_X1 U793 ( .A1(n966), .A2(n702), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n710) );
  NAND2_X1 U795 ( .A1(n718), .A2(G2072), .ZN(n705) );
  NAND2_X1 U796 ( .A1(G1956), .A2(n737), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n519), .A2(n706), .ZN(n711) );
  NOR2_X1 U798 ( .A1(n976), .A2(n711), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U801 ( .A1(n976), .A2(n711), .ZN(n712) );
  XOR2_X1 U802 ( .A(KEYINPUT28), .B(n712), .Z(n713) );
  NOR2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .Z(n717) );
  XNOR2_X1 U805 ( .A(KEYINPUT97), .B(n717), .ZN(n946) );
  NAND2_X1 U806 ( .A1(n718), .A2(n946), .ZN(n719) );
  XNOR2_X1 U807 ( .A(n719), .B(KEYINPUT98), .ZN(n721) );
  INV_X1 U808 ( .A(G1961), .ZN(n1003) );
  NAND2_X1 U809 ( .A1(n1003), .A2(n737), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n729) );
  NAND2_X1 U811 ( .A1(n729), .A2(G171), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n734) );
  NAND2_X1 U813 ( .A1(G8), .A2(n737), .ZN(n810) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n810), .ZN(n724) );
  XOR2_X1 U815 ( .A(KEYINPUT96), .B(n724), .Z(n749) );
  INV_X1 U816 ( .A(G8), .ZN(n725) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n737), .ZN(n748) );
  NOR2_X1 U818 ( .A1(n725), .A2(n748), .ZN(n726) );
  AND2_X1 U819 ( .A1(n749), .A2(n726), .ZN(n727) );
  XOR2_X1 U820 ( .A(n727), .B(KEYINPUT30), .Z(n728) );
  NOR2_X1 U821 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U822 ( .A1(G171), .A2(n729), .ZN(n730) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(n732), .Z(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n736), .B(n735), .ZN(n750) );
  NAND2_X1 U826 ( .A1(n750), .A2(G286), .ZN(n744) );
  NOR2_X1 U827 ( .A1(n737), .A2(G2090), .ZN(n738) );
  XNOR2_X1 U828 ( .A(n738), .B(KEYINPUT104), .ZN(n741) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n810), .ZN(n739) );
  XOR2_X1 U830 ( .A(KEYINPUT103), .B(n739), .Z(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U834 ( .A(KEYINPUT105), .B(n745), .Z(n746) );
  NAND2_X1 U835 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U836 ( .A(n747), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U837 ( .A1(G8), .A2(n748), .ZN(n754) );
  INV_X1 U838 ( .A(n749), .ZN(n752) );
  XOR2_X1 U839 ( .A(n750), .B(KEYINPUT102), .Z(n751) );
  NOR2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n806) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n762), .A2(n757), .ZN(n980) );
  NAND2_X1 U846 ( .A1(n806), .A2(n980), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NOR2_X1 U848 ( .A1(n810), .A2(n758), .ZN(n759) );
  NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n761), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n763), .A2(n810), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n802) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n970) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n824) );
  NAND2_X1 U855 ( .A1(n886), .A2(G128), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G116), .A2(n887), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U858 ( .A(KEYINPUT35), .B(n770), .ZN(n778) );
  XNOR2_X1 U859 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n890), .A2(G104), .ZN(n771) );
  XNOR2_X1 U861 ( .A(n771), .B(KEYINPUT90), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G140), .A2(n859), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT34), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n776), .B(n775), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT36), .B(n779), .Z(n883) );
  XNOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NOR2_X1 U869 ( .A1(n883), .A2(n822), .ZN(n916) );
  NAND2_X1 U870 ( .A1(n824), .A2(n916), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT93), .B(n780), .Z(n820) );
  NAND2_X1 U872 ( .A1(n886), .A2(G119), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G107), .A2(n887), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT94), .B(n783), .Z(n787) );
  NAND2_X1 U876 ( .A1(G95), .A2(n890), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G131), .A2(n859), .ZN(n784) );
  AND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n871) );
  NAND2_X1 U880 ( .A1(G1991), .A2(n871), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G141), .A2(n859), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G129), .A2(n886), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n890), .A2(G105), .ZN(n790) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G117), .A2(n887), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n868) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n868), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n923) );
  NAND2_X1 U891 ( .A1(n923), .A2(n824), .ZN(n797) );
  XNOR2_X1 U892 ( .A(n797), .B(KEYINPUT95), .ZN(n817) );
  INV_X1 U893 ( .A(n817), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n820), .A2(n798), .ZN(n800) );
  XNOR2_X1 U895 ( .A(G1986), .B(G290), .ZN(n982) );
  AND2_X1 U896 ( .A1(n982), .A2(n824), .ZN(n799) );
  NOR2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n803) );
  AND2_X1 U898 ( .A1(n970), .A2(n803), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n829) );
  INV_X1 U900 ( .A(n803), .ZN(n814) );
  NOR2_X1 U901 ( .A1(G2090), .A2(G303), .ZN(n804) );
  NAND2_X1 U902 ( .A1(G8), .A2(n804), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n807), .A2(n810), .ZN(n812) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n808) );
  XOR2_X1 U906 ( .A(n808), .B(KEYINPUT24), .Z(n809) );
  OR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n811) );
  AND2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n827) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n868), .ZN(n931) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n871), .ZN(n919) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n919), .A2(n815), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U915 ( .A1(n931), .A2(n818), .ZN(n819) );
  XNOR2_X1 U916 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n883), .A2(n822), .ZN(n915) );
  NAND2_X1 U919 ( .A1(n823), .A2(n915), .ZN(n825) );
  AND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(n831), .A2(G2106), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n832), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U927 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n838), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U937 ( .A(G261), .ZN(G325) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2072), .B(G2678), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n841), .B(KEYINPUT110), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2100), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1956), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(G1981), .B(G1966), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2474), .B(KEYINPUT111), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(KEYINPUT41), .B(n856), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(n1003), .ZN(G229) );
  NAND2_X1 U959 ( .A1(n887), .A2(G112), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT112), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G100), .A2(n890), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G136), .A2(n859), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n886), .A2(G124), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(n862), .Z(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U968 ( .A(KEYINPUT113), .B(n867), .ZN(G162) );
  XNOR2_X1 U969 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n868), .B(G162), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n874) );
  XNOR2_X1 U972 ( .A(G164), .B(n871), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(n920), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n885) );
  NAND2_X1 U975 ( .A1(n886), .A2(G127), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G115), .A2(n887), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT47), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G139), .A2(n859), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n890), .A2(G103), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n880), .Z(n881) );
  NOR2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n926) );
  XNOR2_X1 U984 ( .A(n883), .B(n926), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n898) );
  NAND2_X1 U986 ( .A1(n886), .A2(G130), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G118), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G106), .A2(n890), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G142), .A2(n859), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n893), .Z(n894) );
  NOR2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U994 ( .A(G160), .B(n896), .Z(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G286), .B(n985), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n904) );
  XOR2_X1 U999 ( .A(n902), .B(G171), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n914), .ZN(n906) );
  XOR2_X1 U1003 ( .A(KEYINPUT115), .B(n906), .Z(n910) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT116), .B(n907), .Z(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT117), .B(n911), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n914), .ZN(G319) );
  INV_X1 U1013 ( .A(n915), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n925) );
  XOR2_X1 U1015 ( .A(G160), .B(G2084), .Z(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n936) );
  XOR2_X1 U1020 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(KEYINPUT50), .B(n929), .ZN(n934) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n932), .Z(n933) );
  NAND2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  INV_X1 U1030 ( .A(KEYINPUT55), .ZN(n962) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n962), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n939), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1033 ( .A(G2090), .B(G35), .Z(n956) );
  XNOR2_X1 U1034 ( .A(G1991), .B(G25), .ZN(n951) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G2072), .B(G33), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(KEYINPUT118), .B(n942), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n943), .B(G32), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G27), .B(n946), .Z(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n949), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(n953), .B(KEYINPUT120), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n954), .B(KEYINPUT53), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(n957), .B(KEYINPUT121), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G2084), .B(G34), .Z(n958) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1054 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n965), .ZN(n1022) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XOR2_X1 U1058 ( .A(G171), .B(G1961), .Z(n968) );
  XNOR2_X1 U1059 ( .A(n966), .B(G1348), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n969), .B(KEYINPUT122), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n973) );
  XOR2_X1 U1064 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n972) );
  XNOR2_X1 U1065 ( .A(n973), .B(n972), .ZN(n984) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G1956), .B(n976), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n985), .ZN(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n1020) );
  INV_X1 U1077 ( .A(G16), .ZN(n1018) );
  XOR2_X1 U1078 ( .A(G1348), .B(KEYINPUT59), .Z(n992) );
  XNOR2_X1 U1079 ( .A(G4), .B(n992), .ZN(n1001) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G20), .ZN(n998) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(KEYINPUT124), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G6), .B(G1981), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(KEYINPUT125), .B(n996), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT126), .B(n999), .Z(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT60), .B(n1002), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1003), .B(G5), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1015) );
  XOR2_X1 U1092 ( .A(G1966), .B(G21), .Z(n1013) );
  XNOR2_X1 U1093 ( .A(G1986), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT127), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT58), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1106 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

