//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n549, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G125), .ZN(new_n459));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(KEYINPUT65), .A2(G113), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n471), .A2(G136), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT66), .ZN(new_n480));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n469), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n476), .B(new_n480), .C1(G124), .C2(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n469), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n469), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n460), .A2(new_n461), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n489), .A2(new_n469), .A3(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(KEYINPUT67), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n487), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n484), .B2(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(G543), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n505), .A2(KEYINPUT68), .A3(G50), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT68), .B1(new_n505), .B2(G50), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT69), .B1(KEYINPUT70), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT69), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n513), .B2(new_n509), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n502), .A2(new_n503), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n516), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n505), .A2(G51), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(G651), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n522), .A2(G90), .B1(G52), .B2(new_n505), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n505), .A2(G43), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n516), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n519), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT73), .ZN(G188));
  AOI22_X1  g127(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n519), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n505), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g135(.A(KEYINPUT74), .B(new_n555), .C1(new_n504), .C2(new_n557), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n516), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT75), .B1(new_n554), .B2(new_n563), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  INV_X1    g144(.A(G166), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n514), .A2(new_n515), .A3(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n505), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n514), .A2(G61), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n575), .A2(new_n576), .B1(G73), .B2(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n514), .A2(KEYINPUT76), .A3(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n522), .A2(G86), .B1(G48), .B2(new_n505), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n519), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n505), .A2(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n516), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n522), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n519), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G54), .B2(new_n505), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n590), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G286), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n568), .B(KEYINPUT77), .Z(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G297));
  AOI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n597), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g185(.A(G2104), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G2105), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n492), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(G2100), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT78), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n484), .A2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n471), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n469), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n616), .B2(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n618), .A2(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2430), .Z(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  AND2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  OAI21_X1  g221(.A(G14), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(KEYINPUT82), .A3(new_n646), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT84), .Z(new_n659));
  INV_X1    g234(.A(new_n657), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n654), .A2(new_n655), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT19), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(KEYINPUT85), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  INV_X1    g262(.A(G34), .ZN(new_n688));
  AOI21_X1  g263(.A(G29), .B1(new_n688), .B2(KEYINPUT24), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(KEYINPUT24), .B2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n473), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G2084), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT96), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(G32), .ZN(new_n696));
  NAND3_X1  g271(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT26), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G129), .B2(new_n484), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n471), .A2(G141), .B1(G105), .B2(new_n612), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(new_n691), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT27), .B(G1996), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G28), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n711), .B1(new_n691), .B2(new_n623), .C1(new_n692), .C2(new_n693), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G1966), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G128), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n471), .A2(G140), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n469), .A2(G116), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n691), .A2(G26), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2067), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n713), .A2(new_n717), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G35), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G162), .B2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n695), .B(new_n730), .C1(new_n731), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n716), .A2(G1966), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT95), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n691), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n691), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT97), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n736), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n546), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1341), .ZN(new_n747));
  NOR2_X1   g322(.A1(G171), .A2(new_n714), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G5), .B2(new_n714), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n747), .B1(G1961), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n691), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n492), .A2(G127), .ZN(new_n753));
  NAND2_X1  g328(.A1(G115), .A2(G2104), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n469), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT25), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n471), .A2(G139), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n755), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(new_n691), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT94), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G2072), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G2072), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n735), .B2(new_n731), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n763), .B(new_n765), .C1(new_n766), .C2(new_n749), .ZN(new_n767));
  NOR2_X1   g342(.A1(G4), .A2(G16), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n597), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT92), .B(G1348), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n769), .B(new_n770), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n714), .A2(G20), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT23), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n568), .B2(new_n714), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1956), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n741), .A2(new_n742), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n771), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n744), .A2(new_n751), .A3(new_n767), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT34), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n780));
  NAND2_X1  g355(.A1(G288), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT90), .A4(new_n573), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G16), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n714), .A2(G23), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT33), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1976), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G22), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G166), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT91), .B(G1971), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n787), .A2(G1976), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(G6), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G305), .B2(new_n714), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT32), .Z(new_n798));
  INV_X1    g373(.A(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n779), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n800), .A2(new_n793), .A3(new_n779), .A4(new_n794), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G24), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n588), .B(KEYINPUT88), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT89), .B(G1986), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G119), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT87), .Z(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G107), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G131), .B2(new_n471), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G25), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n807), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT36), .B1(new_n801), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n800), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n793), .A2(new_n794), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT34), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n824), .A2(new_n825), .A3(new_n802), .A4(new_n819), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n778), .B1(new_n821), .B2(new_n826), .ZN(G311));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n828));
  XNOR2_X1  g403(.A(G311), .B(new_n828), .ZN(G150));
  NAND2_X1  g404(.A1(new_n597), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n519), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT100), .B(G55), .Z(new_n835));
  OAI22_X1  g410(.A1(new_n516), .A2(new_n834), .B1(new_n504), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n546), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n543), .A2(new_n545), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n833), .B2(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n831), .B(new_n841), .Z(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n837), .A2(new_n844), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  INV_X1    g424(.A(G37), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n760), .B(new_n701), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n722), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n500), .A2(KEYINPUT101), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n495), .A2(new_n499), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n814), .B(new_n614), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n484), .A2(G130), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n469), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G142), .B2(new_n471), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n859), .B(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(new_n865), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G160), .B(new_n623), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G162), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n867), .A3(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n874));
  OAI221_X1 g449(.A(new_n850), .B1(new_n868), .B2(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(G299), .B(new_n597), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT103), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n841), .B(new_n607), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n597), .B(new_n568), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n880), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n783), .B(new_n588), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(KEYINPUT104), .ZN(new_n889));
  XNOR2_X1  g464(.A(G305), .B(G303), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(KEYINPUT104), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n887), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n887), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n837), .ZN(G331));
  NAND3_X1  g474(.A1(new_n838), .A2(G301), .A3(new_n840), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G301), .B1(new_n838), .B2(new_n840), .ZN(new_n902));
  OAI21_X1  g477(.A(G286), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G168), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n877), .ZN(new_n907));
  INV_X1    g482(.A(new_n893), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n885), .A2(new_n903), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n850), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n906), .A2(new_n878), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n882), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n881), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n884), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n914), .B(new_n893), .C1(new_n906), .C2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n910), .A4(new_n850), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT44), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n850), .A3(new_n910), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n911), .A2(KEYINPUT43), .A3(new_n912), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n930), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT125), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n814), .A2(new_n817), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n701), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n722), .B(new_n728), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n814), .A2(new_n817), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  AND2_X1   g516(.A1(G290), .A2(G1986), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT45), .B1(new_n857), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n468), .A2(new_n472), .A3(G40), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n468), .A2(new_n472), .A3(KEYINPUT107), .A4(G40), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n943), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(G303), .A2(G8), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT55), .ZN(new_n955));
  INV_X1    g530(.A(G1971), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n500), .A2(new_n944), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n950), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n958), .A2(G1384), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n853), .A2(new_n855), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n956), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(KEYINPUT50), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n495), .B2(new_n499), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n950), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT108), .B(G2090), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n964), .B(KEYINPUT109), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n948), .A2(new_n949), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n958), .B2(new_n957), .ZN(new_n975));
  AOI21_X1  g550(.A(G1971), .B1(new_n975), .B2(new_n962), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n969), .A2(new_n971), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n955), .A2(new_n972), .A3(new_n978), .A4(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n580), .A2(new_n799), .A3(new_n581), .ZN(new_n981));
  INV_X1    g556(.A(new_n581), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n519), .B1(new_n577), .B2(new_n578), .ZN(new_n983));
  OAI21_X1  g558(.A(G1981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT49), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n948), .A2(new_n966), .A3(new_n949), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n981), .B2(new_n984), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n980), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n981), .A2(new_n984), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n986), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(KEYINPUT112), .A3(new_n990), .A4(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  OAI211_X1 g573(.A(G8), .B(new_n989), .C1(new_n783), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n1000));
  INV_X1    g575(.A(G288), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(G1976), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n999), .B2(KEYINPUT52), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n999), .A2(new_n1004), .A3(KEYINPUT52), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n954), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n976), .B2(new_n977), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n979), .A2(new_n997), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT124), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1007), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1016), .A2(new_n1005), .B1(new_n999), .B2(new_n1002), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n993), .B2(new_n996), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT124), .A3(new_n979), .A4(new_n1012), .ZN(new_n1019));
  INV_X1    g594(.A(G1966), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n500), .A2(new_n961), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(new_n960), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n950), .A2(new_n965), .A3(new_n693), .A4(new_n968), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(G168), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1024), .A2(new_n1025), .A3(G8), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(G168), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT51), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(G301), .B(KEYINPUT54), .Z(new_n1032));
  NAND3_X1  g607(.A1(new_n975), .A2(new_n742), .A3(new_n962), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1033), .A2(new_n1034), .B1(new_n766), .B2(new_n969), .ZN(new_n1035));
  OR4_X1    g610(.A1(new_n1034), .A2(new_n960), .A3(G2078), .A4(new_n1021), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n946), .A2(new_n1034), .A3(G2078), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n962), .A2(new_n1038), .ZN(new_n1039));
  OR3_X1    g614(.A1(new_n945), .A2(KEYINPUT123), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT123), .B1(new_n945), .B2(new_n1039), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1032), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n1015), .A2(new_n1019), .A3(new_n1031), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n948), .B(new_n949), .C1(new_n966), .C2(new_n967), .ZN(new_n1046));
  AOI211_X1 g621(.A(KEYINPUT50), .B(G1384), .C1(new_n495), .C2(new_n499), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n770), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n950), .A2(new_n728), .A3(new_n966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT116), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1045), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1045), .A3(new_n1053), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n597), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1056), .B2(new_n597), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1048), .A2(new_n1052), .A3(new_n1049), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1052), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1062), .A3(KEYINPUT60), .ZN(new_n1063));
  INV_X1    g638(.A(new_n597), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT122), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1056), .A2(new_n1057), .A3(new_n597), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1054), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n962), .A2(new_n950), .A3(new_n959), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(new_n564), .B(KEYINPUT57), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n564), .B(KEYINPUT57), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n1072), .A3(new_n1070), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT61), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1075), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT58), .B(G1341), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n989), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT118), .B(G1996), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n962), .A2(new_n950), .A3(new_n959), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n989), .A2(KEYINPUT119), .A3(new_n1083), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n546), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1093), .A3(new_n546), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1092), .A2(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1082), .A2(KEYINPUT121), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT121), .B1(new_n1082), .B2(new_n1097), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1068), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1051), .A2(new_n597), .A3(new_n1053), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1101), .A2(KEYINPUT117), .B1(new_n1074), .B2(new_n1073), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(KEYINPUT117), .B2(new_n1101), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1077), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1044), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1036), .A2(new_n1035), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G286), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(G8), .A3(new_n1024), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1026), .B1(new_n1111), .B2(KEYINPUT51), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1031), .A2(KEYINPUT62), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1015), .A3(new_n1019), .A4(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1117));
  NAND3_X1  g692(.A1(new_n1109), .A2(G8), .A3(G168), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1013), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n972), .A2(new_n978), .A3(G8), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1010), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1018), .A2(new_n1121), .A3(new_n979), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(new_n981), .B(KEYINPUT113), .Z(new_n1126));
  AND2_X1   g701(.A1(new_n993), .A2(new_n996), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1001), .A2(new_n998), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT114), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n979), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1130), .A2(new_n990), .B1(new_n1018), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1116), .A2(new_n1125), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n953), .B1(new_n1106), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n951), .A2(new_n935), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT46), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n937), .A2(new_n702), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n952), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT47), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n951), .A2(new_n940), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n951), .A2(new_n941), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT48), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n722), .A2(G2067), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n938), .B2(new_n933), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n952), .A2(new_n1147), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1140), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n932), .B1(new_n1134), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1140), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1116), .A2(new_n1125), .A3(new_n1132), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1099), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1082), .A2(KEYINPUT121), .A3(new_n1097), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1104), .B1(new_n1155), .B2(new_n1068), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1152), .B1(new_n1156), .B2(new_n1044), .ZN(new_n1157));
  OAI211_X1 g732(.A(KEYINPUT125), .B(new_n1151), .C1(new_n1157), .C2(new_n953), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1150), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n1161));
  NOR2_X1   g735(.A1(G227), .A2(new_n457), .ZN(new_n1162));
  XOR2_X1   g736(.A(new_n1162), .B(KEYINPUT126), .Z(new_n1163));
  OR3_X1    g737(.A1(G401), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g738(.A(new_n1161), .B1(G401), .B2(new_n1163), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n875), .A2(new_n686), .ZN(new_n1167));
  INV_X1    g741(.A(new_n1167), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n1166), .A2(new_n922), .A3(new_n1168), .ZN(G308));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n922), .A3(new_n1168), .ZN(G225));
endmodule


