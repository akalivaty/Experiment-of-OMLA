//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  OR2_X1    g000(.A1(KEYINPUT66), .A2(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT66), .A2(G119), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G116), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n187), .A2(new_n190), .A3(G116), .A4(new_n188), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n196), .A3(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT65), .A2(G131), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G131), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(new_n206), .A3(new_n207), .A4(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n207), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n205), .A2(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n215), .A3(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT1), .B1(new_n220), .B2(G146), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n218), .A2(new_n219), .B1(G128), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n210), .B(new_n213), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n210), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT64), .B1(new_n220), .B2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n220), .A2(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n219), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n233), .A2(new_n236), .B1(new_n234), .B2(new_n223), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n227), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n227), .B2(new_n238), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n200), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n227), .A2(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(new_n199), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n196), .B1(new_n193), .B2(new_n194), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n242), .A2(new_n247), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT31), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n243), .A2(KEYINPUT28), .A3(new_n246), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n227), .A2(new_n238), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n200), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT28), .B1(new_n243), .B2(new_n246), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n242), .A2(new_n263), .A3(new_n247), .A4(new_n254), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G472), .A2(G902), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(KEYINPUT69), .A3(new_n266), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(KEYINPUT32), .A3(new_n266), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n265), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n266), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n279));
  INV_X1    g093(.A(new_n261), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n259), .A3(new_n257), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n281), .B2(new_n253), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n242), .A2(new_n247), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n254), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n278), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n246), .A2(KEYINPUT70), .A3(new_n238), .A4(new_n227), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n259), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT70), .B1(new_n243), .B2(new_n246), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND4_X1   g104(.A1(KEYINPUT29), .A2(new_n290), .A3(new_n280), .A4(new_n254), .ZN(new_n291));
  OAI21_X1  g105(.A(G472), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n272), .A2(new_n277), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G137), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(G221), .A3(G234), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n294), .B(new_n296), .Z(new_n297));
  AND2_X1   g111(.A1(KEYINPUT66), .A2(G119), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT66), .A2(G119), .ZN(new_n299));
  OAI21_X1  g113(.A(G128), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G119), .A2(G128), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(KEYINPUT23), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G110), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n224), .B1(new_n298), .B2(new_n299), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT24), .B(G110), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n300), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  INV_X1    g127(.A(G125), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT16), .ZN(new_n316));
  OR3_X1    g130(.A1(new_n314), .A2(KEYINPUT16), .A3(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G146), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n215), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n309), .B1(new_n300), .B2(new_n302), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n215), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n326), .B2(new_n318), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n303), .A2(new_n307), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G110), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n297), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n332));
  INV_X1    g146(.A(new_n309), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n224), .B1(new_n187), .B2(new_n188), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n301), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n316), .A2(G146), .A3(new_n317), .ZN(new_n336));
  AOI21_X1  g150(.A(G146), .B1(new_n316), .B2(new_n317), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n304), .B1(new_n303), .B2(new_n307), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n321), .B1(new_n308), .B2(new_n310), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n323), .A2(new_n330), .A3(KEYINPUT73), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n331), .B1(new_n344), .B2(new_n297), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G234), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n347), .B2(G217), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(KEYINPUT25), .C1(new_n345), .C2(G902), .ZN(new_n351));
  OAI21_X1  g165(.A(G217), .B1(new_n347), .B2(G902), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT72), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n297), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n342), .B2(new_n343), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n278), .B1(new_n356), .B2(new_n331), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT25), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n349), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n293), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G140), .ZN(new_n362));
  INV_X1    g176(.A(G227), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G953), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n362), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n368));
  AOI21_X1  g182(.A(G101), .B1(new_n367), .B2(G107), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G104), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n367), .A2(G107), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n366), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n221), .A2(G128), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n233), .A2(new_n379), .B1(new_n223), .B2(new_n225), .ZN(new_n380));
  INV_X1    g194(.A(new_n377), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT77), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n223), .B1(G128), .B2(new_n221), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n382), .B(new_n381), .C1(new_n385), .C2(new_n226), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n384), .A2(KEYINPUT78), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT78), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  INV_X1    g202(.A(new_n230), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT79), .B1(new_n390), .B2(KEYINPUT12), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n386), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT78), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n230), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT79), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT12), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n389), .A2(new_n398), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n391), .A2(new_n399), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n368), .A2(new_n372), .A3(new_n376), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G101), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT4), .A3(new_n382), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n405), .A2(new_n237), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n386), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT10), .B1(new_n222), .B2(new_n226), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n378), .A2(new_n383), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n408), .A2(new_n414), .A3(new_n230), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n365), .B1(new_n401), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n408), .A2(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n389), .ZN(new_n418));
  INV_X1    g232(.A(new_n365), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n230), .B1(new_n408), .B2(new_n414), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n416), .A2(G469), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n391), .A2(new_n399), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n392), .A2(new_n400), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n419), .B1(new_n418), .B2(new_n421), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n426), .B(new_n278), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G469), .A2(G902), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n425), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G214), .B1(G237), .B2(G902), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n434), .B(KEYINPUT80), .Z(new_n435));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n193), .B2(new_n194), .ZN(new_n438));
  OAI21_X1  g252(.A(G113), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n198), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n440), .B2(new_n413), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(KEYINPUT81), .A3(new_n198), .A4(new_n412), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n405), .A2(new_n200), .A3(new_n407), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n441), .A2(new_n443), .A3(new_n446), .A4(new_n444), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n380), .A2(new_n314), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n314), .B2(new_n237), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT82), .B(G224), .Z(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n295), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT83), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n454), .B(new_n457), .Z(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(new_n454), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n440), .B1(new_n373), .B2(new_n377), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n413), .B2(new_n440), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n446), .B(KEYINPUT8), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n465), .B2(new_n449), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n459), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n435), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G237), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n295), .A3(G214), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(new_n220), .ZN(new_n476));
  AOI21_X1  g290(.A(G143), .B1(new_n249), .B2(G214), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT18), .A2(G131), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n313), .A2(new_n315), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G146), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n478), .A2(new_n479), .B1(new_n320), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n220), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n479), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT85), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n488), .B(new_n479), .C1(new_n483), .C2(new_n484), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n482), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n203), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n476), .B2(new_n477), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n203), .A3(new_n484), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n480), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n319), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n496), .B(new_n215), .C1(new_n498), .C2(new_n495), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n499), .A3(new_n318), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n490), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n490), .A2(new_n500), .A3(KEYINPUT87), .ZN(new_n504));
  XOR2_X1   g318(.A(G113), .B(G122), .Z(new_n505));
  XOR2_X1   g319(.A(KEYINPUT88), .B(G104), .Z(new_n506));
  XOR2_X1   g320(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n492), .A2(new_n511), .A3(new_n493), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n485), .A2(KEYINPUT17), .A3(new_n491), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n326), .A3(new_n318), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n490), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n510), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n514), .A2(new_n490), .A3(KEYINPUT89), .A4(new_n507), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n503), .A2(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT90), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n503), .A2(new_n508), .A3(new_n504), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n522), .A3(new_n519), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n515), .A2(new_n508), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n278), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n533), .A2(G475), .B1(new_n526), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n220), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n224), .A2(G143), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n205), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n191), .A2(G122), .ZN(new_n540));
  INV_X1    g354(.A(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G116), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n542), .A3(new_n371), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n371), .B1(new_n540), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n220), .A2(KEYINPUT13), .A3(G128), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(new_n538), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n537), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n205), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT14), .B1(new_n541), .B2(G116), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n541), .A2(G116), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT91), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n191), .B2(G122), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n540), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n557), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G107), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n537), .A2(new_n538), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G134), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n544), .B1(new_n565), .B2(new_n539), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n563), .A2(KEYINPUT92), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT92), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n553), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n347), .A2(KEYINPUT9), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n347), .A2(KEYINPUT9), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT9), .B(G234), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT75), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n295), .A2(G217), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT93), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT93), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT94), .B1(new_n569), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n558), .A2(new_n540), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n585), .A2(KEYINPUT91), .B1(new_n557), .B2(new_n555), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n371), .B1(new_n586), .B2(new_n560), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n565), .A2(new_n539), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n543), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n563), .A2(KEYINPUT92), .A3(new_n566), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n552), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n581), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n569), .A2(new_n582), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n278), .ZN(new_n597));
  INV_X1    g411(.A(G478), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(KEYINPUT15), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n295), .A2(G952), .ZN(new_n601));
  NAND2_X1  g415(.A1(G234), .A2(G237), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT21), .B(G898), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT95), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(G902), .A3(G953), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT96), .Z(new_n608));
  OAI211_X1 g422(.A(new_n596), .B(new_n278), .C1(KEYINPUT15), .C2(new_n598), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n600), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n536), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n573), .A2(new_n575), .A3(new_n278), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G221), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n433), .A2(new_n473), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n361), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n374), .ZN(G3));
  NAND2_X1  g430(.A1(new_n265), .A2(new_n278), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G472), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n269), .A2(new_n618), .A3(new_n271), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n359), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(new_n613), .A3(new_n433), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n581), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n579), .A2(KEYINPUT97), .A3(new_n580), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT98), .B1(new_n592), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n592), .B2(new_n581), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n569), .A2(new_n629), .A3(new_n623), .A4(new_n624), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT99), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n626), .A2(new_n628), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n596), .A2(new_n627), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n598), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT100), .B1(new_n597), .B2(new_n598), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n597), .A2(KEYINPUT100), .A3(new_n598), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n638), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n536), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n467), .A2(new_n468), .ZN(new_n644));
  INV_X1    g458(.A(new_n435), .ZN(new_n645));
  INV_X1    g459(.A(new_n468), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n459), .A2(new_n466), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n608), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n621), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND2_X1  g467(.A1(new_n600), .A2(new_n609), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n533), .A2(G475), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n534), .A2(new_n522), .ZN(new_n656));
  INV_X1    g470(.A(new_n529), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n648), .A2(new_n658), .A3(new_n649), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n621), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(new_n344), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n297), .A2(KEYINPUT36), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n348), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n354), .B2(new_n358), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n619), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n614), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT37), .B(G110), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NAND2_X1  g488(.A1(new_n293), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n433), .A2(new_n613), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n675), .A2(new_n676), .A3(new_n648), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n602), .A2(new_n678), .A3(G902), .A4(G953), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT101), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT101), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n603), .A3(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n655), .B(new_n682), .C1(new_n657), .C2(new_n656), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n600), .B2(new_n609), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  INV_X1    g500(.A(new_n676), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n682), .B(KEYINPUT39), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n459), .A2(new_n471), .A3(new_n466), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n471), .B1(new_n459), .B2(new_n466), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n693), .B(new_n694), .Z(new_n695));
  AND2_X1   g509(.A1(new_n272), .A2(new_n277), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n253), .B1(new_n288), .B2(new_n289), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n255), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n698), .B2(KEYINPUT103), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(KEYINPUT103), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G472), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n536), .A2(new_n654), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n435), .A3(new_n668), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n695), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n690), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NAND3_X1  g522(.A1(new_n642), .A2(new_n536), .A3(new_n682), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n677), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  AND2_X1   g526(.A1(new_n293), .A2(new_n360), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n428), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n420), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n430), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(G469), .B1(new_n718), .B2(G902), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(new_n613), .A3(new_n431), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n713), .A2(new_n650), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NAND3_X1  g537(.A1(new_n713), .A2(new_n659), .A3(new_n720), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  INV_X1    g540(.A(new_n648), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n726), .B1(new_n720), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n613), .A3(new_n431), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n648), .A3(KEYINPUT104), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n293), .A2(new_n668), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n611), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(G119), .Z(G21));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n256), .A2(new_n264), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n254), .B1(new_n290), .B2(new_n280), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n266), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT106), .B(G472), .Z(new_n740));
  AOI22_X1  g554(.A1(new_n736), .A2(new_n739), .B1(new_n617), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(KEYINPUT105), .B(new_n266), .C1(new_n737), .C2(new_n738), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n360), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n360), .A2(new_n741), .A3(new_n745), .A4(new_n742), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n648), .A2(new_n703), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n729), .A2(new_n649), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n736), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n617), .A2(new_n740), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n668), .A2(new_n752), .A3(new_n742), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n741), .A2(KEYINPUT108), .A3(new_n668), .A4(new_n742), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n709), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n728), .B2(new_n730), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  NOR3_X1   g574(.A1(new_n691), .A2(new_n692), .A3(new_n435), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n293), .A2(new_n360), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n676), .A2(KEYINPUT109), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n433), .A2(new_n764), .A3(new_n613), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT42), .B1(new_n766), .B2(new_n710), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n267), .A2(new_n270), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n292), .A2(new_n273), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT42), .A3(new_n360), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n709), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n433), .A2(new_n764), .A3(new_n613), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n764), .B1(new_n433), .B2(new_n613), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n771), .B(new_n761), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n293), .A2(new_n360), .A3(new_n761), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n710), .C1(new_n773), .C2(new_n772), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n774), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  OAI211_X1 g598(.A(new_n777), .B(new_n684), .C1(new_n773), .C2(new_n772), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n419), .B1(new_n716), .B2(new_n418), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n423), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n416), .A2(KEYINPUT45), .A3(new_n424), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n790), .A3(G469), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n432), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(KEYINPUT46), .A3(new_n432), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n431), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n613), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(new_n688), .ZN(new_n799));
  INV_X1    g613(.A(new_n639), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n632), .A2(new_n634), .B1(new_n627), .B2(new_n596), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n800), .A2(new_n640), .B1(new_n801), .B2(new_n637), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT43), .B1(new_n802), .B2(new_n536), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT43), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n530), .A2(new_n535), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n642), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n619), .A2(new_n668), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n761), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT44), .B1(new_n807), .B2(new_n808), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n799), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  NOR2_X1   g630(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n797), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n796), .B(new_n613), .C1(new_n820), .C2(new_n817), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n709), .A2(new_n812), .A3(new_n293), .A4(new_n360), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  NOR2_X1   g638(.A1(G952), .A2(G953), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n683), .A2(new_n654), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n433), .A2(new_n761), .A3(new_n827), .A4(new_n613), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n675), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n766), .B2(new_n684), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n758), .B(new_n761), .C1(new_n773), .C2(new_n772), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT114), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n829), .ZN(new_n833));
  AND4_X1   g647(.A1(KEYINPUT114), .A2(new_n785), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n776), .B(new_n782), .C1(new_n832), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT112), .B1(new_n642), .B2(new_n536), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n654), .A2(new_n530), .A3(new_n535), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n802), .B2(new_n805), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(KEYINPUT112), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n645), .B(new_n608), .C1(new_n691), .C2(new_n692), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n620), .A3(new_n613), .A4(new_n433), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n614), .B1(new_n361), .B2(new_n671), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT113), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n643), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n654), .A2(new_n530), .A3(new_n535), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n536), .B2(new_n642), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n849), .B2(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n621), .A3(new_n841), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  INV_X1    g666(.A(new_n614), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n713), .B2(new_n670), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n727), .A2(new_n433), .A3(new_n613), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n857), .B(new_n732), .C1(new_n684), .C2(new_n710), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n682), .B(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n669), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n687), .A2(new_n702), .A3(new_n748), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n759), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n750), .A2(new_n721), .A3(new_n724), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n734), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n858), .A2(new_n759), .A3(new_n867), .A4(new_n862), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n856), .A2(new_n864), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n826), .B1(new_n835), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n868), .A2(new_n856), .A3(new_n864), .A4(new_n866), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT53), .B1(new_n767), .B2(new_n775), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n785), .A2(new_n831), .A3(new_n833), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n830), .A2(KEYINPUT114), .A3(new_n831), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n876), .A2(new_n877), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n783), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n871), .B1(new_n882), .B2(new_n870), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n720), .A2(new_n761), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n702), .A2(new_n885), .A3(new_n359), .A4(new_n603), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n536), .A3(new_n642), .ZN(new_n887));
  INV_X1    g701(.A(new_n603), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n803), .A2(new_n888), .A3(new_n806), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n803), .A2(new_n891), .A3(new_n806), .A4(new_n888), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n890), .A2(new_n892), .B1(new_n746), .B2(new_n744), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n887), .B(new_n601), .C1(new_n894), .C2(new_n731), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n885), .B1(new_n890), .B2(new_n892), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n769), .A2(new_n360), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n898), .A2(KEYINPUT48), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(KEYINPUT48), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n719), .A2(new_n431), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n613), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n819), .B2(new_n821), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n893), .A2(new_n761), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT51), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n756), .A2(new_n757), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n642), .A2(new_n536), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n896), .A2(new_n907), .B1(new_n886), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n695), .A2(new_n645), .A3(new_n729), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n893), .A2(KEYINPUT50), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT50), .B1(new_n893), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n901), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n904), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n918));
  INV_X1    g732(.A(new_n905), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT117), .B1(new_n904), .B2(new_n905), .ZN(new_n921));
  OAI211_X1 g735(.A(KEYINPUT118), .B(new_n909), .C1(new_n911), .C2(new_n912), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n916), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n914), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n825), .B1(new_n884), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n360), .A2(new_n613), .A3(new_n645), .ZN(new_n927));
  OR4_X1    g741(.A1(new_n536), .A2(new_n695), .A3(new_n802), .A4(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n902), .B(KEYINPUT49), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n702), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT119), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n882), .A2(new_n870), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n925), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n825), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  INV_X1    g752(.A(new_n930), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n931), .A2(new_n940), .ZN(G75));
  NOR2_X1   g755(.A1(new_n295), .A2(G952), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n278), .B1(new_n870), .B2(new_n879), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT56), .B1(new_n944), .B2(G210), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n450), .A2(new_n452), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n458), .ZN(new_n947));
  XNOR2_X1  g761(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n945), .B2(new_n950), .ZN(G51));
  NAND2_X1  g766(.A1(new_n870), .A2(new_n879), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n934), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n432), .B(KEYINPUT57), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n430), .B2(new_n429), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n791), .B(KEYINPUT121), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n944), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n942), .B1(new_n958), .B2(new_n960), .ZN(G54));
  AND3_X1   g775(.A1(new_n944), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n943), .B1(new_n962), .B2(new_n528), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n528), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT122), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n962), .A2(new_n966), .A3(new_n528), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n963), .B1(new_n965), .B2(new_n967), .ZN(G60));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT59), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n955), .A2(new_n801), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n933), .A2(new_n934), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n801), .B1(new_n972), .B2(new_n970), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n971), .A2(new_n973), .A3(new_n942), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n870), .B2(new_n879), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n665), .A3(new_n666), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n978), .B(new_n943), .C1(new_n346), .C2(new_n977), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G66));
  AOI21_X1  g795(.A(new_n295), .B1(new_n605), .B2(new_n455), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n856), .A2(new_n866), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n295), .ZN(new_n984));
  INV_X1    g798(.A(G898), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n946), .B1(new_n985), .B2(G953), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G69));
  OAI21_X1  g801(.A(G953), .B1(new_n363), .B2(new_n678), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n798), .A2(new_n688), .A3(new_n748), .A4(new_n897), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n858), .A2(new_n759), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(new_n785), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n815), .A2(new_n990), .A3(new_n823), .A4(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n783), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n295), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n678), .A2(G953), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n240), .A2(new_n241), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n496), .B1(new_n498), .B2(new_n495), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT123), .Z(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n995), .A2(new_n996), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n689), .A2(new_n839), .A3(new_n762), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n799), .B2(new_n814), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n707), .A2(new_n991), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n707), .A2(new_n1007), .A3(new_n991), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1004), .A2(new_n1006), .A3(new_n823), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1000), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n295), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1001), .A2(new_n1002), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1002), .B1(new_n1001), .B2(new_n1011), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n989), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1014), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n988), .A3(new_n1012), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(G72));
  NOR2_X1   g832(.A1(new_n283), .A2(new_n254), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n993), .A2(new_n994), .A3(new_n983), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1019), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1022), .B1(new_n1009), .B2(new_n983), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT125), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n284), .A2(new_n253), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1024), .B(new_n943), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1027), .A2(new_n1023), .A3(new_n1019), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n932), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1032), .A2(KEYINPUT126), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(KEYINPUT126), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(G57));
endmodule


