//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  AOI21_X1  g050(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(G136), .ZN(new_n478));
  MUX2_X1   g053(.A(G100), .B(G112), .S(G2105), .Z(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  MUX2_X1   g057(.A(G102), .B(G114), .S(G2105), .Z(new_n483));
  AOI22_X1  g058(.A1(G126), .A2(new_n476), .B1(new_n483), .B2(G2104), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n467), .A2(new_n485), .A3(G138), .ZN(new_n486));
  INV_X1    g061(.A(new_n466), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n461), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT67), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n467), .A2(new_n493), .A3(G138), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n491), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI211_X1 g070(.A(KEYINPUT68), .B(new_n493), .C1(new_n486), .C2(new_n490), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n484), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n502), .A2(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n514), .B(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n511), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n510), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n508), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n499), .B2(new_n500), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(G89), .B1(G51), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n505), .A2(new_n504), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n525), .A2(new_n526), .A3(G63), .A4(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n527), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G90), .Z(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n519), .A2(new_n533), .B1(G52), .B2(new_n521), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n525), .A2(new_n526), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G651), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n535), .B1(new_n545), .B2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n502), .A2(new_n548), .B1(new_n508), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n537), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(KEYINPUT74), .A3(G651), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n521), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n523), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(G651), .A2(new_n569), .B1(new_n519), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n545), .A2(new_n546), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(new_n534), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n537), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n519), .A2(G87), .B1(G49), .B2(new_n521), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n521), .A2(G48), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n508), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n511), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n519), .A2(G85), .B1(G47), .B2(new_n521), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n525), .A2(new_n526), .A3(G60), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT76), .B1(new_n591), .B2(G651), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  AOI211_X1 g168(.A(new_n593), .B(new_n511), .C1(new_n589), .C2(new_n590), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n588), .B1(new_n592), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n508), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n501), .A2(new_n512), .A3(KEYINPUT10), .A4(G92), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(G66), .B1(new_n505), .B2(new_n504), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n602), .A2(KEYINPUT77), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT77), .B1(new_n602), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n602), .A2(new_n606), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n602), .A2(KEYINPUT77), .A3(new_n606), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n612), .A2(KEYINPUT78), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n596), .B1(G868), .B2(new_n615), .ZN(G284));
  XNOR2_X1  g191(.A(G284), .B(KEYINPUT79), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  MUX2_X1   g193(.A(G286), .B(G299), .S(new_n618), .Z(G297));
  MUX2_X1   g194(.A(G286), .B(G299), .S(new_n618), .Z(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n621), .B2(G860), .ZN(G148));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n615), .B2(new_n621), .ZN(new_n624));
  AOI211_X1 g199(.A(KEYINPUT80), .B(G559), .C1(new_n609), .C2(new_n614), .ZN(new_n625));
  OAI21_X1  g200(.A(G868), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n467), .A2(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  MUX2_X1   g209(.A(G99), .B(G111), .S(G2105), .Z(new_n635));
  AOI22_X1  g210(.A1(G123), .A2(new_n476), .B1(new_n635), .B2(G2104), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n468), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n650), .B2(new_n652), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n647), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n666), .B2(new_n660), .ZN(new_n667));
  INV_X1    g242(.A(new_n660), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n667), .B1(new_n668), .B2(new_n665), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n660), .A2(new_n661), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n659), .B1(new_n670), .B2(KEYINPUT17), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n664), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n639), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n632), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  AOI211_X1 g259(.A(new_n682), .B(new_n684), .C1(new_n677), .C2(new_n681), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G23), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n579), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G6), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n586), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n697), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT85), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G290), .B2(new_n693), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  MUX2_X1   g291(.A(G95), .B(G107), .S(G2105), .Z(new_n717));
  AOI22_X1  g292(.A1(G119), .A2(new_n476), .B1(new_n717), .B2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(G131), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n468), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT83), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n721), .B(new_n723), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n715), .A2(new_n716), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n707), .B2(new_n708), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n711), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n728), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n711), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n693), .A2(G20), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT23), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G299), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1956), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  AOI22_X1  g314(.A1(G128), .A2(new_n476), .B1(new_n467), .B2(G140), .ZN(new_n740));
  MUX2_X1   g315(.A(G104), .B(G116), .S(G2105), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2104), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(KEYINPUT89), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(KEYINPUT89), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT90), .B(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n737), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT93), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G160), .B2(G29), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G2084), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n638), .A2(new_n737), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT31), .B(G11), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT96), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT30), .B(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n737), .B2(new_n758), .ZN(new_n759));
  AND4_X1   g334(.A1(new_n748), .A2(new_n754), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n753), .A2(G2084), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT27), .B(G1996), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n737), .A2(G32), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT26), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n467), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n476), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(G29), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n761), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n760), .B(new_n772), .C1(new_n763), .C2(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G16), .B2(G21), .ZN(new_n776));
  NOR2_X1   g351(.A1(G286), .A2(new_n693), .ZN(new_n777));
  MUX2_X1   g352(.A(new_n776), .B(new_n775), .S(new_n777), .Z(new_n778));
  AOI211_X1 g353(.A(new_n736), .B(new_n773), .C1(new_n774), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n615), .B2(G16), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1348), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n467), .A2(G139), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT25), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(KEYINPUT25), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT91), .Z(new_n788));
  AOI22_X1  g363(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n461), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G33), .B(new_n792), .S(G29), .Z(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G2072), .Z(new_n794));
  NAND3_X1  g369(.A1(new_n779), .A2(new_n782), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n778), .A2(new_n774), .ZN(new_n796));
  NOR2_X1   g371(.A1(G29), .A2(G35), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G162), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT29), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n796), .B1(G2090), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G2090), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(G164), .A2(G29), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G27), .B2(G29), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(G2078), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G5), .A2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G301), .B2(new_n693), .ZN(new_n808));
  INV_X1    g383(.A(G1961), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n803), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n805), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G16), .A2(G19), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n558), .B2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT88), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1341), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n781), .A2(G1348), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n795), .A2(new_n814), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n729), .A2(new_n731), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND3_X1  g397(.A1(new_n525), .A2(new_n526), .A3(G67), .ZN(new_n823));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n511), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n502), .A2(new_n826), .B1(new_n508), .B2(new_n827), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n825), .A2(KEYINPUT98), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT98), .B1(new_n825), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  INV_X1    g408(.A(new_n558), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n834), .A2(KEYINPUT99), .A3(new_n830), .A4(new_n829), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n825), .A2(new_n828), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n558), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n558), .A2(new_n831), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n615), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(G860), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n833), .B1(new_n849), .B2(new_n850), .ZN(G145));
  XNOR2_X1  g426(.A(KEYINPUT103), .B(G37), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n497), .A2(KEYINPUT101), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n493), .B1(new_n486), .B2(new_n490), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n494), .A2(new_n492), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n484), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n745), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n630), .B(new_n720), .ZN(new_n864));
  MUX2_X1   g439(.A(G106), .B(G118), .S(G2105), .Z(new_n865));
  AOI22_X1  g440(.A1(G130), .A2(new_n476), .B1(new_n865), .B2(G2104), .ZN(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n468), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n864), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n863), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n792), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n770), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n869), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n863), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n854), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G160), .B(new_n481), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(new_n638), .Z(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n853), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n874), .A2(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n881), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT40), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n883), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G395));
  XOR2_X1   g464(.A(G299), .B(new_n610), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n624), .B2(new_n625), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n607), .A2(new_n608), .A3(new_n597), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT78), .B1(new_n612), .B2(new_n613), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n621), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT80), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n615), .A2(new_n623), .A3(new_n621), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(KEYINPUT105), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n893), .A2(new_n899), .A3(new_n840), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n840), .B1(new_n893), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n838), .A2(new_n839), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n558), .A2(new_n831), .A3(new_n836), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n624), .A2(new_n625), .A3(new_n892), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT105), .B1(new_n897), .B2(new_n898), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n893), .A2(new_n899), .A3(new_n840), .ZN(new_n909));
  INV_X1    g484(.A(new_n890), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(G288), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n579), .B(new_n588), .C1(new_n592), .C2(new_n594), .ZN(new_n913));
  XNOR2_X1  g488(.A(G303), .B(new_n586), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n913), .ZN(new_n920));
  INV_X1    g495(.A(new_n914), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(KEYINPUT42), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n902), .A2(new_n911), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n902), .B2(new_n911), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI211_X1 g506(.A(KEYINPUT107), .B(new_n927), .C1(new_n902), .C2(new_n911), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n831), .A2(new_n618), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g511(.A1(G295), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(KEYINPUT108), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  INV_X1    g515(.A(new_n923), .ZN(new_n941));
  NAND2_X1  g516(.A1(G301), .A2(G286), .ZN(new_n942));
  NAND2_X1  g517(.A1(G171), .A2(G168), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n840), .ZN(new_n944));
  NOR2_X1   g519(.A1(G171), .A2(G168), .ZN(new_n945));
  AOI211_X1 g520(.A(G286), .B(new_n535), .C1(new_n545), .C2(new_n546), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n905), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n947), .A3(new_n890), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n891), .B1(new_n944), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n941), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n944), .A2(new_n947), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n923), .B(new_n948), .C1(new_n953), .C2(new_n891), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n954), .A3(new_n852), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n954), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n940), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n957), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n951), .A2(new_n954), .A3(KEYINPUT43), .A4(new_n958), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n862), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G160), .A2(G40), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n745), .B(G2067), .Z(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n770), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(KEYINPUT109), .A3(new_n974), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n720), .A2(new_n723), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n720), .A2(new_n723), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(G290), .B(G1986), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n970), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT120), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n497), .A2(new_n986), .A3(KEYINPUT45), .A4(new_n965), .ZN(new_n987));
  INV_X1    g562(.A(new_n969), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n859), .B2(new_n484), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n987), .B(new_n988), .C1(KEYINPUT45), .C2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n986), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n774), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n497), .A2(new_n965), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n969), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n497), .A2(new_n995), .A3(new_n965), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT116), .B(G2084), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n994), .A2(new_n997), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n985), .B(G8), .C1(new_n1002), .C2(G286), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G168), .A2(G8), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n992), .B2(new_n1001), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G168), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n985), .B(new_n1005), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n969), .B1(new_n993), .B2(new_n967), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n855), .A2(KEYINPUT45), .A3(new_n861), .A4(new_n965), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1971), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n988), .B1(new_n989), .B2(new_n995), .ZN(new_n1016));
  INV_X1    g591(.A(new_n996), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(new_n1017), .A3(G2090), .ZN(new_n1018));
  OAI21_X1  g593(.A(G8), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(new_n1021), .C2(new_n1020), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n994), .A2(new_n997), .A3(new_n999), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(G8), .B(new_n1025), .C1(new_n1030), .C2(new_n1015), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(G1981), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n586), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(G1981), .B1(new_n583), .B2(new_n585), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT49), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n497), .A2(new_n965), .A3(new_n988), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n579), .A2(G1976), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n579), .B2(G1976), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1037), .A2(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT112), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1041), .A2(new_n1047), .A3(KEYINPUT52), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1044), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1027), .A2(new_n1031), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n994), .A2(new_n999), .A3(new_n997), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT122), .B(G1961), .Z(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT123), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT123), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1061));
  NOR2_X1   g636(.A1(G171), .A2(new_n1061), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n969), .B(KEYINPUT124), .Z(new_n1064));
  NAND2_X1  g639(.A1(new_n968), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT125), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n968), .A2(new_n1067), .A3(new_n1064), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1052), .A2(G2078), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1066), .A2(new_n1014), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1063), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n990), .A2(new_n991), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1072), .A2(new_n1069), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1054), .ZN(new_n1074));
  OR2_X1    g649(.A1(G301), .A2(new_n1061), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n1075), .C1(KEYINPUT54), .C2(G171), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1012), .A2(new_n1051), .A3(new_n1071), .A4(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1038), .A2(G2067), .ZN(new_n1078));
  INV_X1    g653(.A(G1348), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1055), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n607), .A2(new_n608), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1080), .B2(KEYINPUT60), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n735), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1013), .A2(new_n1014), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(G299), .B(KEYINPUT57), .Z(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1013), .A2(new_n1014), .A3(new_n972), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n1038), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1096), .B1(new_n1100), .B2(new_n558), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT59), .B(new_n834), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1095), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1086), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1094), .A2(KEYINPUT118), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1087), .A2(new_n1089), .A3(new_n1106), .A4(new_n1091), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT61), .B1(new_n1108), .B2(new_n1093), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(KEYINPUT119), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1111), .B(KEYINPUT61), .C1(new_n1108), .C2(new_n1093), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1104), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1093), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1108), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1077), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT114), .Z(new_n1118));
  NOR2_X1   g693(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1033), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(G8), .A3(new_n1038), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1049), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1031), .ZN(new_n1123));
  AND4_X1   g698(.A1(KEYINPUT63), .A2(new_n1031), .A3(new_n1007), .A4(new_n1049), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1053), .A2(new_n704), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1029), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1127), .B2(G8), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT117), .B(new_n1008), .C1(new_n1126), .C2(new_n1029), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1026), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1007), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1050), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1123), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1004), .A2(new_n1137), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1074), .A2(G171), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1050), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1135), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n984), .B1(new_n1116), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n982), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n982), .A2(new_n1144), .ZN(new_n1146));
  NOR4_X1   g721(.A1(new_n968), .A2(G1986), .A3(G290), .A4(new_n969), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT48), .Z(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n980), .B(KEYINPUT126), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n977), .A2(new_n978), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n745), .A2(G2067), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n970), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n971), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n970), .B1(new_n770), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT46), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n970), .B2(new_n972), .ZN(new_n1157));
  NOR4_X1   g732(.A1(new_n968), .A2(KEYINPUT46), .A3(G1996), .A4(new_n969), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1149), .A2(new_n1153), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1143), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g737(.A1(G401), .A2(new_n459), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n691), .A2(new_n674), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g739(.A(new_n1165), .B1(new_n883), .B2(new_n886), .ZN(new_n1166));
  NAND3_X1  g740(.A1(new_n1166), .A2(new_n961), .A3(new_n962), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


