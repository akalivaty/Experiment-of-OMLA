

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(n528), .B(n527), .ZN(n874) );
  XNOR2_X1 U553 ( .A(n524), .B(n523), .ZN(n526) );
  NOR2_X1 U554 ( .A1(n799), .A2(n747), .ZN(n520) );
  BUF_X1 U555 ( .A(n714), .Z(n725) );
  NOR2_X1 U556 ( .A1(G1966), .A2(n799), .ZN(n736) );
  XNOR2_X1 U557 ( .A(n522), .B(KEYINPUT23), .ZN(n523) );
  AND2_X1 U558 ( .A1(n521), .A2(G2104), .ZN(n873) );
  NOR2_X1 U559 ( .A1(G651), .A2(n617), .ZN(n638) );
  XOR2_X1 U560 ( .A(KEYINPUT65), .B(n533), .Z(G160) );
  INV_X1 U561 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U562 ( .A1(G101), .A2(n873), .ZN(n524) );
  INV_X1 U563 ( .A(KEYINPUT66), .ZN(n522) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n521), .ZN(n870) );
  NAND2_X1 U565 ( .A1(G125), .A2(n870), .ZN(n525) );
  NAND2_X1 U566 ( .A1(n526), .A2(n525), .ZN(n532) );
  XNOR2_X1 U567 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n528) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  NAND2_X1 U569 ( .A1(G137), .A2(n874), .ZN(n530) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U571 ( .A1(G113), .A2(n871), .ZN(n529) );
  NAND2_X1 U572 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U573 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U575 ( .A1(n642), .A2(G89), .ZN(n534) );
  XNOR2_X1 U576 ( .A(n534), .B(KEYINPUT4), .ZN(n536) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n617) );
  INV_X1 U578 ( .A(G651), .ZN(n538) );
  NOR2_X1 U579 ( .A1(n617), .A2(n538), .ZN(n640) );
  NAND2_X1 U580 ( .A1(G76), .A2(n640), .ZN(n535) );
  NAND2_X1 U581 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U582 ( .A(n537), .B(KEYINPUT5), .ZN(n545) );
  NAND2_X1 U583 ( .A1(n638), .A2(G51), .ZN(n542) );
  NOR2_X1 U584 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U585 ( .A(KEYINPUT68), .B(n539), .Z(n540) );
  XNOR2_X1 U586 ( .A(KEYINPUT1), .B(n540), .ZN(n645) );
  NAND2_X1 U587 ( .A1(G63), .A2(n645), .ZN(n541) );
  NAND2_X1 U588 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U589 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U590 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U591 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U593 ( .A1(n638), .A2(G52), .ZN(n548) );
  NAND2_X1 U594 ( .A1(G64), .A2(n645), .ZN(n547) );
  NAND2_X1 U595 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U596 ( .A1(G90), .A2(n642), .ZN(n550) );
  NAND2_X1 U597 ( .A1(G77), .A2(n640), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U600 ( .A1(n553), .A2(n552), .ZN(G171) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G108), .ZN(G238) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  NAND2_X1 U606 ( .A1(G94), .A2(G452), .ZN(n554) );
  XOR2_X1 U607 ( .A(KEYINPUT70), .B(n554), .Z(G173) );
  NAND2_X1 U608 ( .A1(G7), .A2(G661), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U610 ( .A(G223), .ZN(n823) );
  NAND2_X1 U611 ( .A1(n823), .A2(G567), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT73), .ZN(n557) );
  XNOR2_X1 U613 ( .A(KEYINPUT11), .B(n557), .ZN(G234) );
  NAND2_X1 U614 ( .A1(n642), .A2(G81), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G68), .A2(n640), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U618 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n561) );
  XNOR2_X1 U619 ( .A(n562), .B(n561), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G56), .A2(n645), .ZN(n563) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n563), .Z(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n638), .A2(G43), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n928) );
  INV_X1 U625 ( .A(G860), .ZN(n607) );
  OR2_X1 U626 ( .A1(n928), .A2(n607), .ZN(G153) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G54), .A2(n638), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n642), .A2(G92), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G66), .A2(n645), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G79), .A2(n640), .ZN(n570) );
  XNOR2_X1 U633 ( .A(KEYINPUT75), .B(n570), .ZN(n571) );
  NOR2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U636 ( .A(n575), .B(KEYINPUT15), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT76), .B(n576), .Z(n849) );
  NOR2_X1 U638 ( .A1(n849), .A2(G868), .ZN(n578) );
  INV_X1 U639 ( .A(G868), .ZN(n659) );
  NOR2_X1 U640 ( .A1(n659), .A2(G301), .ZN(n577) );
  NOR2_X1 U641 ( .A1(n578), .A2(n577), .ZN(G284) );
  NAND2_X1 U642 ( .A1(G78), .A2(n640), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n642), .A2(G91), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G65), .A2(n645), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G53), .A2(n638), .ZN(n581) );
  XNOR2_X1 U647 ( .A(KEYINPUT71), .B(n581), .ZN(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT72), .ZN(G299) );
  NOR2_X1 U651 ( .A1(G286), .A2(n659), .ZN(n588) );
  NOR2_X1 U652 ( .A1(G299), .A2(G868), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(G297) );
  NAND2_X1 U654 ( .A1(n607), .A2(G559), .ZN(n589) );
  INV_X1 U655 ( .A(n849), .ZN(n919) );
  NAND2_X1 U656 ( .A1(n589), .A2(n919), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n590), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U658 ( .A1(G868), .A2(n928), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n919), .A2(G868), .ZN(n591) );
  NOR2_X1 U660 ( .A1(G559), .A2(n591), .ZN(n592) );
  NOR2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G282) );
  XOR2_X1 U662 ( .A(G2100), .B(KEYINPUT80), .Z(n605) );
  NAND2_X1 U663 ( .A1(G123), .A2(n870), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT18), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G135), .A2(n874), .ZN(n595) );
  XOR2_X1 U666 ( .A(KEYINPUT77), .B(n595), .Z(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n873), .A2(G99), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT78), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G111), .A2(n871), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT79), .B(n601), .Z(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n992) );
  XNOR2_X1 U674 ( .A(n992), .B(G2096), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U676 ( .A1(n919), .A2(G559), .ZN(n606) );
  XOR2_X1 U677 ( .A(n928), .B(n606), .Z(n656) );
  NAND2_X1 U678 ( .A1(n607), .A2(n656), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n640), .A2(G80), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G67), .A2(n645), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G93), .A2(n642), .ZN(n610) );
  XNOR2_X1 U683 ( .A(KEYINPUT81), .B(n610), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n638), .A2(G55), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n658) );
  XNOR2_X1 U687 ( .A(n615), .B(n658), .ZN(G145) );
  NAND2_X1 U688 ( .A1(G74), .A2(G651), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(KEYINPUT82), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G49), .A2(n638), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G87), .A2(n617), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n645), .A2(n620), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U695 ( .A1(G50), .A2(n638), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n640), .A2(G75), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G62), .A2(n645), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G88), .A2(n642), .ZN(n625) );
  XNOR2_X1 U700 ( .A(KEYINPUT85), .B(n625), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n630), .B(KEYINPUT86), .ZN(G303) );
  NAND2_X1 U704 ( .A1(G85), .A2(n642), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G72), .A2(n640), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U707 ( .A1(G60), .A2(n645), .ZN(n633) );
  XNOR2_X1 U708 ( .A(KEYINPUT69), .B(n633), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(G47), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U712 ( .A1(G48), .A2(n638), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n639), .B(KEYINPUT84), .ZN(n650) );
  NAND2_X1 U714 ( .A1(G73), .A2(n640), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n642), .A2(G86), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U718 ( .A1(G61), .A2(n645), .ZN(n646) );
  XNOR2_X1 U719 ( .A(KEYINPUT83), .B(n646), .ZN(n647) );
  NOR2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U722 ( .A(G288), .B(KEYINPUT19), .ZN(n652) );
  XNOR2_X1 U723 ( .A(G299), .B(G303), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(G290), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(n658), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(G305), .ZN(n848) );
  XNOR2_X1 U728 ( .A(n656), .B(n848), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U738 ( .A1(G236), .A2(G238), .ZN(n666) );
  NAND2_X1 U739 ( .A1(G69), .A2(n666), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n667), .A2(G237), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT87), .ZN(n828) );
  NAND2_X1 U742 ( .A1(G567), .A2(n828), .ZN(n673) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U745 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G96), .A2(n671), .ZN(n827) );
  NAND2_X1 U747 ( .A1(G2106), .A2(n827), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT88), .B(n674), .Z(G319) );
  INV_X1 U750 ( .A(G319), .ZN(n676) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U752 ( .A1(n676), .A2(n675), .ZN(n826) );
  NAND2_X1 U753 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(n874), .A2(G138), .ZN(n679) );
  NAND2_X1 U755 ( .A1(G102), .A2(n873), .ZN(n677) );
  XOR2_X1 U756 ( .A(KEYINPUT89), .B(n677), .Z(n678) );
  NAND2_X1 U757 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U758 ( .A1(G114), .A2(n871), .ZN(n681) );
  NAND2_X1 U759 ( .A1(G126), .A2(n870), .ZN(n680) );
  NAND2_X1 U760 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U761 ( .A1(n683), .A2(n682), .ZN(G164) );
  NOR2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n921) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n750) );
  AND2_X1 U764 ( .A1(G40), .A2(n750), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G160), .A2(n684), .ZN(n685) );
  XNOR2_X2 U766 ( .A(n685), .B(KEYINPUT64), .ZN(n714) );
  INV_X1 U767 ( .A(n714), .ZN(n709) );
  NAND2_X1 U768 ( .A1(G2067), .A2(n709), .ZN(n687) );
  NAND2_X1 U769 ( .A1(n714), .A2(G1348), .ZN(n686) );
  NAND2_X1 U770 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U771 ( .A(n688), .B(KEYINPUT99), .ZN(n695) );
  OR2_X1 U772 ( .A1(n919), .A2(n695), .ZN(n694) );
  XOR2_X1 U773 ( .A(G1996), .B(KEYINPUT98), .Z(n943) );
  NOR2_X1 U774 ( .A1(n714), .A2(n943), .ZN(n689) );
  XOR2_X1 U775 ( .A(n689), .B(KEYINPUT26), .Z(n691) );
  NAND2_X1 U776 ( .A1(n725), .A2(G1341), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n928), .A2(n692), .ZN(n693) );
  NAND2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U780 ( .A1(n919), .A2(n695), .ZN(n696) );
  NAND2_X1 U781 ( .A1(n697), .A2(n696), .ZN(n703) );
  INV_X1 U782 ( .A(KEYINPUT27), .ZN(n699) );
  NAND2_X1 U783 ( .A1(G2072), .A2(n709), .ZN(n698) );
  XNOR2_X1 U784 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U785 ( .A1(n725), .A2(G1956), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U787 ( .A1(G299), .A2(n704), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U789 ( .A1(G299), .A2(n704), .ZN(n705) );
  XOR2_X1 U790 ( .A(KEYINPUT28), .B(n705), .Z(n706) );
  NOR2_X1 U791 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U792 ( .A(n708), .B(KEYINPUT29), .ZN(n713) );
  XNOR2_X1 U793 ( .A(KEYINPUT25), .B(G2078), .ZN(n952) );
  NAND2_X1 U794 ( .A1(n709), .A2(n952), .ZN(n711) );
  XNOR2_X1 U795 ( .A(G1961), .B(KEYINPUT97), .ZN(n964) );
  NAND2_X1 U796 ( .A1(n725), .A2(n964), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n711), .A2(n710), .ZN(n718) );
  NAND2_X1 U798 ( .A1(G171), .A2(n718), .ZN(n712) );
  NAND2_X1 U799 ( .A1(n713), .A2(n712), .ZN(n723) );
  NAND2_X1 U800 ( .A1(n714), .A2(G8), .ZN(n799) );
  NOR2_X1 U801 ( .A1(n725), .A2(G2084), .ZN(n733) );
  NOR2_X1 U802 ( .A1(n736), .A2(n733), .ZN(n715) );
  NAND2_X1 U803 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U804 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U805 ( .A1(G168), .A2(n717), .ZN(n720) );
  NOR2_X1 U806 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U808 ( .A(KEYINPUT31), .B(n721), .Z(n722) );
  NAND2_X1 U809 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U810 ( .A(n724), .B(KEYINPUT100), .ZN(n734) );
  NAND2_X1 U811 ( .A1(n734), .A2(G286), .ZN(n730) );
  NOR2_X1 U812 ( .A1(n725), .A2(G2090), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n799), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n728), .A2(G303), .ZN(n729) );
  NAND2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U817 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U818 ( .A(n732), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U819 ( .A1(G8), .A2(n733), .ZN(n738) );
  INV_X1 U820 ( .A(n734), .ZN(n735) );
  NOR2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U823 ( .A1(n740), .A2(n739), .ZN(n793) );
  NOR2_X1 U824 ( .A1(G303), .A2(G1971), .ZN(n741) );
  XNOR2_X1 U825 ( .A(KEYINPUT101), .B(n741), .ZN(n742) );
  NAND2_X1 U826 ( .A1(n793), .A2(n742), .ZN(n743) );
  NOR2_X1 U827 ( .A1(n921), .A2(n743), .ZN(n745) );
  NAND2_X1 U828 ( .A1(G288), .A2(G1976), .ZN(n744) );
  XOR2_X1 U829 ( .A(KEYINPUT102), .B(n744), .Z(n920) );
  NOR2_X1 U830 ( .A1(n745), .A2(n920), .ZN(n746) );
  XNOR2_X1 U831 ( .A(n746), .B(KEYINPUT103), .ZN(n786) );
  XOR2_X1 U832 ( .A(G1981), .B(G305), .Z(n924) );
  INV_X1 U833 ( .A(n924), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n921), .A2(KEYINPUT33), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n748), .A2(n520), .ZN(n783) );
  NAND2_X1 U836 ( .A1(G160), .A2(G40), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n816) );
  NAND2_X1 U838 ( .A1(G104), .A2(n873), .ZN(n752) );
  NAND2_X1 U839 ( .A1(G140), .A2(n874), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U841 ( .A(KEYINPUT34), .B(n753), .ZN(n759) );
  NAND2_X1 U842 ( .A1(G116), .A2(n871), .ZN(n755) );
  NAND2_X1 U843 ( .A1(G128), .A2(n870), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U845 ( .A(KEYINPUT35), .B(n756), .Z(n757) );
  XNOR2_X1 U846 ( .A(KEYINPUT90), .B(n757), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U848 ( .A(KEYINPUT36), .B(n760), .ZN(n897) );
  XNOR2_X1 U849 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  OR2_X1 U850 ( .A1(n897), .A2(n814), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n761), .B(KEYINPUT91), .ZN(n1013) );
  NAND2_X1 U852 ( .A1(n816), .A2(n1013), .ZN(n812) );
  NAND2_X1 U853 ( .A1(G107), .A2(n871), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G119), .A2(n870), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U856 ( .A(KEYINPUT92), .B(n764), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G95), .A2(n873), .ZN(n766) );
  NAND2_X1 U858 ( .A1(G131), .A2(n874), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n885) );
  INV_X1 U861 ( .A(G1991), .ZN(n804) );
  NOR2_X1 U862 ( .A1(n885), .A2(n804), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G141), .A2(n874), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G129), .A2(n870), .ZN(n769) );
  NAND2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U866 ( .A1(G105), .A2(n873), .ZN(n771) );
  XNOR2_X1 U867 ( .A(n771), .B(KEYINPUT93), .ZN(n772) );
  XNOR2_X1 U868 ( .A(n772), .B(KEYINPUT38), .ZN(n773) );
  NOR2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n871), .A2(G117), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n888) );
  AND2_X1 U872 ( .A1(G1996), .A2(n888), .ZN(n777) );
  NOR2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n994) );
  XOR2_X1 U874 ( .A(n816), .B(KEYINPUT94), .Z(n779) );
  NOR2_X1 U875 ( .A1(n994), .A2(n779), .ZN(n809) );
  XNOR2_X1 U876 ( .A(KEYINPUT95), .B(n809), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n812), .A2(n780), .ZN(n782) );
  XNOR2_X1 U878 ( .A(G1986), .B(G290), .ZN(n938) );
  AND2_X1 U879 ( .A1(n938), .A2(n816), .ZN(n781) );
  NOR2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n790) );
  AND2_X1 U881 ( .A1(n783), .A2(n790), .ZN(n787) );
  INV_X1 U882 ( .A(n787), .ZN(n784) );
  OR2_X1 U883 ( .A1(n799), .A2(n784), .ZN(n785) );
  NOR2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n789) );
  AND2_X1 U885 ( .A1(n787), .A2(KEYINPUT33), .ZN(n788) );
  NOR2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n821) );
  INV_X1 U887 ( .A(n790), .ZN(n803) );
  NOR2_X1 U888 ( .A1(G303), .A2(G2090), .ZN(n791) );
  NAND2_X1 U889 ( .A1(G8), .A2(n791), .ZN(n792) );
  XNOR2_X1 U890 ( .A(n792), .B(KEYINPUT104), .ZN(n794) );
  NAND2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n795) );
  AND2_X1 U892 ( .A1(n795), .A2(n799), .ZN(n801) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U894 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  XNOR2_X1 U895 ( .A(KEYINPUT96), .B(n797), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n819) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n888), .ZN(n998) );
  AND2_X1 U900 ( .A1(n804), .A2(n885), .ZN(n996) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n805) );
  XOR2_X1 U902 ( .A(n805), .B(KEYINPUT105), .Z(n806) );
  NOR2_X1 U903 ( .A1(n996), .A2(n806), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT106), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n998), .A2(n810), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n814), .A2(n897), .ZN(n1000) );
  NAND2_X1 U910 ( .A1(n815), .A2(n1000), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U917 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(G188) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT108), .ZN(G325) );
  XNOR2_X1 U923 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  XOR2_X1 U925 ( .A(G2100), .B(KEYINPUT43), .Z(n831) );
  XNOR2_X1 U926 ( .A(G2090), .B(G2678), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U928 ( .A(n832), .B(KEYINPUT42), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U931 ( .A(KEYINPUT110), .B(G2096), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1976), .B(G1981), .Z(n840) );
  XNOR2_X1 U936 ( .A(G1966), .B(G1961), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U938 ( .A(n841), .B(G2474), .Z(n843) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1956), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U941 ( .A(KEYINPUT41), .B(G1971), .Z(n845) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U945 ( .A(n848), .B(G286), .Z(n851) );
  XNOR2_X1 U946 ( .A(G171), .B(n849), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n852), .B(n928), .ZN(n853) );
  NOR2_X1 U949 ( .A1(G37), .A2(n853), .ZN(G397) );
  NAND2_X1 U950 ( .A1(G124), .A2(n870), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n873), .A2(G100), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G136), .A2(n874), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G112), .A2(n871), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U957 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U958 ( .A1(n871), .A2(G115), .ZN(n861) );
  XOR2_X1 U959 ( .A(KEYINPUT115), .B(n861), .Z(n863) );
  NAND2_X1 U960 ( .A1(n870), .A2(G127), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT47), .B(n864), .ZN(n869) );
  NAND2_X1 U963 ( .A1(G103), .A2(n873), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G139), .A2(n874), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U966 ( .A(KEYINPUT114), .B(n867), .Z(n868) );
  NAND2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n1002) );
  NAND2_X1 U968 ( .A1(G130), .A2(n870), .ZN(n882) );
  NAND2_X1 U969 ( .A1(n871), .A2(G118), .ZN(n872) );
  XNOR2_X1 U970 ( .A(KEYINPUT111), .B(n872), .ZN(n880) );
  NAND2_X1 U971 ( .A1(G106), .A2(n873), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U974 ( .A(KEYINPUT112), .B(n877), .Z(n878) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n878), .ZN(n879) );
  NOR2_X1 U976 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n883), .B(n992), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n1002), .B(n884), .ZN(n887) );
  XNOR2_X1 U980 ( .A(G160), .B(n885), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n887), .B(n886), .ZN(n891) );
  XOR2_X1 U982 ( .A(G164), .B(n888), .Z(n889) );
  XNOR2_X1 U983 ( .A(n889), .B(G162), .ZN(n890) );
  XOR2_X1 U984 ( .A(n891), .B(n890), .Z(n896) );
  XOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n893) );
  XNOR2_X1 U986 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U988 ( .A(KEYINPUT116), .B(n894), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U991 ( .A1(G37), .A2(n899), .ZN(n900) );
  XNOR2_X1 U992 ( .A(KEYINPUT118), .B(n900), .ZN(G395) );
  XOR2_X1 U993 ( .A(KEYINPUT107), .B(G2451), .Z(n902) );
  XNOR2_X1 U994 ( .A(G2446), .B(G2427), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(n909) );
  XOR2_X1 U996 ( .A(G2438), .B(G2435), .Z(n904) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2430), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(n905), .B(G2454), .Z(n907) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(n910), .A2(G14), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(n917), .A2(G319), .ZN(n914) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n912), .B(KEYINPUT119), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G397), .A2(G395), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  INV_X1 U1013 ( .A(n917), .ZN(G401) );
  INV_X1 U1014 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U1015 ( .A(G16), .B(KEYINPUT124), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(KEYINPUT56), .ZN(n942) );
  XNOR2_X1 U1017 ( .A(G1348), .B(n919), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n934) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G168), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(n926), .B(KEYINPUT125), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT57), .B(n927), .Z(n932) );
  XNOR2_X1 U1024 ( .A(n928), .B(G1341), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(G299), .B(G1956), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n940) );
  XNOR2_X1 U1029 ( .A(G171), .B(G1961), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(G166), .B(G1971), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n1023) );
  XNOR2_X1 U1035 ( .A(n943), .B(G32), .ZN(n951) );
  XNOR2_X1 U1036 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(G25), .B(G1991), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(G28), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(KEYINPUT122), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(G33), .B(n947), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G27), .B(n952), .Z(n953) );
  NOR2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1046 ( .A(KEYINPUT53), .B(n955), .Z(n959) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(G34), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n956), .B(KEYINPUT123), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G2084), .B(n957), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n987) );
  NAND2_X1 U1053 ( .A1(KEYINPUT55), .A2(n987), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n962), .ZN(n1021) );
  XOR2_X1 U1055 ( .A(G5), .B(KEYINPUT126), .Z(n963) );
  XNOR2_X1 U1056 ( .A(n964), .B(n963), .ZN(n971) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1060 ( .A(G1986), .B(G24), .Z(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT58), .B(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n982) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(KEYINPUT59), .B(G4), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n972), .B(KEYINPUT127), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(G1348), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G20), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G6), .B(G1981), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT60), .B(n980), .Z(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G21), .B(G1966), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n985), .Z(n986) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n986), .ZN(n990) );
  OR2_X1 U1079 ( .A1(KEYINPUT55), .A2(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1019) );
  XOR2_X1 U1082 ( .A(G160), .B(G2084), .Z(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1011) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n999), .Z(n1001) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1009) );
  XNOR2_X1 U1090 ( .A(KEYINPUT120), .B(n1002), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(G2072), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(G164), .B(G2078), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT121), .B(n1006), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1014), .ZN(n1016) );
  INV_X1 U1100 ( .A(KEYINPUT55), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(G29), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1105 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

