

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U322 ( .A(n397), .B(n396), .ZN(n404) );
  XNOR2_X1 U323 ( .A(n452), .B(n451), .ZN(n516) );
  XNOR2_X1 U324 ( .A(n475), .B(n474), .ZN(n476) );
  AND2_X1 U325 ( .A1(n444), .A2(n565), .ZN(n420) );
  XNOR2_X1 U326 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n457) );
  XNOR2_X1 U327 ( .A(n458), .B(n457), .ZN(n459) );
  NOR2_X1 U328 ( .A1(n441), .A2(n517), .ZN(n442) );
  INV_X1 U329 ( .A(G197GAT), .ZN(n394) );
  INV_X1 U330 ( .A(KEYINPUT54), .ZN(n470) );
  XNOR2_X1 U331 ( .A(n395), .B(n394), .ZN(n397) );
  XNOR2_X1 U332 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U333 ( .A(n408), .B(n323), .ZN(n409) );
  XNOR2_X1 U334 ( .A(KEYINPUT37), .B(KEYINPUT109), .ZN(n451) );
  XNOR2_X1 U335 ( .A(n410), .B(n409), .ZN(n415) );
  XNOR2_X1 U336 ( .A(n477), .B(n476), .ZN(n561) );
  XNOR2_X1 U337 ( .A(KEYINPUT26), .B(n419), .ZN(n565) );
  XNOR2_X1 U338 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U339 ( .A(n454), .B(G29GAT), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n485), .B(n484), .ZN(G1349GAT) );
  XNOR2_X1 U341 ( .A(n456), .B(n455), .ZN(G1328GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n291) );
  XOR2_X1 U343 ( .A(G141GAT), .B(G22GAT), .Z(n407) );
  XOR2_X1 U344 ( .A(G169GAT), .B(G8GAT), .Z(n383) );
  XNOR2_X1 U345 ( .A(n407), .B(n383), .ZN(n290) );
  XNOR2_X1 U346 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U347 ( .A(n292), .B(G197GAT), .Z(n298) );
  XNOR2_X1 U348 ( .A(G15GAT), .B(G1GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n293), .B(KEYINPUT72), .ZN(n352) );
  XOR2_X1 U350 ( .A(n352), .B(KEYINPUT68), .Z(n295) );
  NAND2_X1 U351 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n296), .B(G113GAT), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n308) );
  XOR2_X1 U355 ( .A(G43GAT), .B(G29GAT), .Z(n300) );
  XNOR2_X1 U356 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U358 ( .A(n301), .B(KEYINPUT71), .Z(n303) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n336) );
  XOR2_X1 U361 ( .A(KEYINPUT73), .B(KEYINPUT30), .Z(n305) );
  XNOR2_X1 U362 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U364 ( .A(n336), .B(n306), .Z(n307) );
  XOR2_X1 U365 ( .A(n308), .B(n307), .Z(n567) );
  XOR2_X1 U366 ( .A(KEYINPUT74), .B(n567), .Z(n532) );
  XOR2_X1 U367 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n310) );
  XNOR2_X1 U368 ( .A(KEYINPUT79), .B(KEYINPUT31), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U370 ( .A(G148GAT), .B(G78GAT), .Z(n402) );
  XOR2_X1 U371 ( .A(KEYINPUT33), .B(n402), .Z(n312) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G71GAT), .Z(n360) );
  XNOR2_X1 U373 ( .A(n360), .B(G204GAT), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U375 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n318) );
  XNOR2_X1 U378 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n317), .B(KEYINPUT75), .ZN(n351) );
  XOR2_X1 U380 ( .A(n318), .B(n351), .Z(n325) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(G64GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n319), .B(KEYINPUT78), .ZN(n386) );
  INV_X1 U383 ( .A(G106GAT), .ZN(n323) );
  XOR2_X1 U384 ( .A(KEYINPUT77), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n386), .B(n329), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n571) );
  NAND2_X1 U390 ( .A1(n532), .A2(n571), .ZN(n492) );
  XNOR2_X1 U391 ( .A(KEYINPUT36), .B(KEYINPUT108), .ZN(n339) );
  XOR2_X1 U392 ( .A(G190GAT), .B(KEYINPUT81), .Z(n389) );
  XOR2_X1 U393 ( .A(KEYINPUT11), .B(KEYINPUT82), .Z(n326) );
  XNOR2_X1 U394 ( .A(n389), .B(n326), .ZN(n327) );
  XOR2_X1 U395 ( .A(G218GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U396 ( .A(n327), .B(n403), .ZN(n328) );
  XOR2_X1 U397 ( .A(n328), .B(KEYINPUT80), .Z(n331) );
  XNOR2_X1 U398 ( .A(G134GAT), .B(n329), .ZN(n330) );
  XNOR2_X1 U399 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U400 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n333) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U402 ( .A(n333), .B(n332), .Z(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n336), .B(KEYINPUT10), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n554) );
  XNOR2_X1 U406 ( .A(KEYINPUT83), .B(n554), .ZN(n486) );
  XNOR2_X1 U407 ( .A(n339), .B(n486), .ZN(n580) );
  XOR2_X1 U408 ( .A(G64GAT), .B(G155GAT), .Z(n341) );
  XNOR2_X1 U409 ( .A(G22GAT), .B(G8GAT), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n356) );
  XOR2_X1 U411 ( .A(G183GAT), .B(KEYINPUT84), .Z(n388) );
  XOR2_X1 U412 ( .A(G78GAT), .B(G211GAT), .Z(n343) );
  XNOR2_X1 U413 ( .A(G127GAT), .B(G71GAT), .ZN(n342) );
  XNOR2_X1 U414 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U415 ( .A(n388), .B(n344), .Z(n346) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U417 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U418 ( .A(KEYINPUT85), .B(KEYINPUT15), .Z(n348) );
  XNOR2_X1 U419 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U421 ( .A(n350), .B(n349), .Z(n354) );
  XNOR2_X1 U422 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U424 ( .A(n356), .B(n355), .Z(n557) );
  XOR2_X1 U425 ( .A(G176GAT), .B(G190GAT), .Z(n358) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(G99GAT), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U428 ( .A(n360), .B(n359), .Z(n362) );
  NAND2_X1 U429 ( .A1(G227GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n364) );
  XNOR2_X1 U432 ( .A(G15GAT), .B(KEYINPUT88), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U434 ( .A(KEYINPUT87), .B(G183GAT), .Z(n366) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(KEYINPUT90), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U437 ( .A(n368), .B(n367), .Z(n374) );
  XOR2_X1 U438 ( .A(G127GAT), .B(KEYINPUT0), .Z(n370) );
  XNOR2_X1 U439 ( .A(G113GAT), .B(G134GAT), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n432) );
  XOR2_X1 U441 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n372) );
  XNOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n371) );
  XNOR2_X1 U443 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n432), .B(n377), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U446 ( .A(n376), .B(n375), .Z(n478) );
  XOR2_X1 U447 ( .A(n377), .B(KEYINPUT97), .Z(n379) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U449 ( .A(n379), .B(n378), .ZN(n393) );
  XOR2_X1 U450 ( .A(KEYINPUT98), .B(KEYINPUT95), .Z(n381) );
  XNOR2_X1 U451 ( .A(G218GAT), .B(G92GAT), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U453 ( .A(n382), .B(KEYINPUT96), .Z(n385) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(n383), .ZN(n384) );
  XNOR2_X1 U455 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U456 ( .A(n387), .B(n386), .Z(n391) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n399) );
  XNOR2_X1 U460 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n395) );
  XOR2_X1 U461 ( .A(KEYINPUT92), .B(G211GAT), .Z(n396) );
  INV_X1 U462 ( .A(n404), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n469) );
  NOR2_X1 U464 ( .A1(n478), .A2(n469), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n400), .B(KEYINPUT101), .ZN(n416) );
  XNOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n401), .B(KEYINPUT2), .ZN(n431) );
  XOR2_X1 U468 ( .A(n431), .B(n402), .Z(n406) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n410) );
  XNOR2_X1 U471 ( .A(G50GAT), .B(n407), .ZN(n408) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n412) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U475 ( .A(KEYINPUT23), .B(n413), .Z(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n473) );
  NAND2_X1 U477 ( .A1(n416), .A2(n473), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n417), .B(KEYINPUT102), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n418), .B(KEYINPUT25), .ZN(n422) );
  INV_X1 U480 ( .A(n469), .ZN(n519) );
  XNOR2_X1 U481 ( .A(KEYINPUT27), .B(n519), .ZN(n444) );
  INV_X1 U482 ( .A(n478), .ZN(n559) );
  NOR2_X1 U483 ( .A1(n559), .A2(n473), .ZN(n419) );
  XNOR2_X1 U484 ( .A(KEYINPUT100), .B(n420), .ZN(n421) );
  NOR2_X1 U485 ( .A1(n422), .A2(n421), .ZN(n441) );
  XOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n424) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(G57GAT), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n440) );
  XOR2_X1 U489 ( .A(G148GAT), .B(G120GAT), .Z(n426) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(G141GAT), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U492 ( .A(G162GAT), .B(G85GAT), .Z(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n436) );
  XNOR2_X1 U494 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n429), .B(KEYINPUT94), .ZN(n430) );
  XOR2_X1 U496 ( .A(n430), .B(KEYINPUT5), .Z(n434) );
  XNOR2_X1 U497 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n438) );
  NAND2_X1 U500 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n517) );
  XNOR2_X1 U503 ( .A(n442), .B(KEYINPUT103), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n443) );
  XNOR2_X1 U505 ( .A(n473), .B(n443), .ZN(n531) );
  NAND2_X1 U506 ( .A1(n517), .A2(n444), .ZN(n528) );
  NOR2_X1 U507 ( .A1(n531), .A2(n528), .ZN(n445) );
  XOR2_X1 U508 ( .A(KEYINPUT99), .B(n445), .Z(n446) );
  NAND2_X1 U509 ( .A1(n446), .A2(n478), .ZN(n447) );
  NAND2_X1 U510 ( .A1(n448), .A2(n447), .ZN(n449) );
  XOR2_X1 U511 ( .A(KEYINPUT104), .B(n449), .Z(n490) );
  NOR2_X1 U512 ( .A1(n557), .A2(n490), .ZN(n450) );
  NAND2_X1 U513 ( .A1(n580), .A2(n450), .ZN(n452) );
  NOR2_X1 U514 ( .A1(n492), .A2(n516), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n453), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U516 ( .A1(n503), .A2(n517), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT110), .B(KEYINPUT39), .Z(n454) );
  NAND2_X1 U518 ( .A1(n580), .A2(n557), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n459), .A2(n571), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT114), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n461), .A2(n532), .ZN(n467) );
  XOR2_X1 U522 ( .A(n571), .B(KEYINPUT41), .Z(n547) );
  NOR2_X1 U523 ( .A1(n567), .A2(n547), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT46), .ZN(n463) );
  NOR2_X1 U525 ( .A1(n557), .A2(n463), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n554), .A2(n464), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U529 ( .A(KEYINPUT48), .B(n468), .ZN(n529) );
  NOR2_X1 U530 ( .A1(n529), .A2(n469), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n517), .A2(n472), .ZN(n566) );
  NAND2_X1 U532 ( .A1(n566), .A2(n473), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n475) );
  INV_X1 U534 ( .A(KEYINPUT55), .ZN(n474) );
  NOR2_X1 U535 ( .A1(n561), .A2(n478), .ZN(n556) );
  NAND2_X1 U536 ( .A1(n556), .A2(n532), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(G169GAT), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1348GAT) );
  INV_X1 U540 ( .A(n547), .ZN(n535) );
  NAND2_X1 U541 ( .A1(n556), .A2(n535), .ZN(n485) );
  XOR2_X1 U542 ( .A(G176GAT), .B(KEYINPUT56), .Z(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n482) );
  INV_X1 U544 ( .A(n557), .ZN(n575) );
  NOR2_X1 U545 ( .A1(n486), .A2(n575), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT86), .B(n487), .Z(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT16), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT105), .B(n491), .ZN(n507) );
  NOR2_X1 U550 ( .A1(n492), .A2(n507), .ZN(n500) );
  NAND2_X1 U551 ( .A1(n517), .A2(n500), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT34), .ZN(n494) );
  XOR2_X1 U553 ( .A(n494), .B(KEYINPUT107), .Z(n496) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(KEYINPUT106), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U556 ( .A1(n500), .A2(n519), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U559 ( .A1(n500), .A2(n559), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n531), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U563 ( .A1(n519), .A2(n503), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n559), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT40), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n503), .A2(n531), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  NAND2_X1 U571 ( .A1(n567), .A2(n535), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n507), .A2(n515), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n512), .A2(n517), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n519), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n559), .A2(n512), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U580 ( .A1(n512), .A2(n531), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U586 ( .A1(n524), .A2(n519), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n559), .A2(n524), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(KEYINPUT112), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n526) );
  NAND2_X1 U592 ( .A1(n524), .A2(n531), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT115), .Z(n534) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n545), .A2(n559), .ZN(n530) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n541), .A2(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U602 ( .A1(n541), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U605 ( .A1(n541), .A2(n557), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U609 ( .A1(n541), .A2(n486), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n544), .Z(G1343GAT) );
  NAND2_X1 U612 ( .A1(n545), .A2(n565), .ZN(n553) );
  NOR2_X1 U613 ( .A1(n567), .A2(n553), .ZN(n546) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U615 ( .A1(n547), .A2(n553), .ZN(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n575), .A2(n553), .ZN(n551) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(n551), .Z(n552) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n563) );
  NAND2_X1 U627 ( .A1(n559), .A2(n486), .ZN(n560) );
  OR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(G190GAT), .B(n564), .Z(G1351GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n578) );
  NOR2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n578), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(n576), .Z(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

