//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G169gat), .B(G197gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT12), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT91), .ZN(new_n217));
  INV_X1    g016(.A(G43gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G43gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT15), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT90), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n220), .B2(G43gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n226), .A2(new_n227), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n217), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(new_n222), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G1gat), .B2(new_n233), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g038(.A1(KEYINPUT92), .A2(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT92), .A2(KEYINPUT17), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n232), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n229), .A2(new_n231), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n239), .B1(new_n245), .B2(new_n238), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT93), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT18), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n210), .B1(new_n249), .B2(KEYINPUT97), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n238), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n236), .B(G8gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT95), .B1(new_n257), .B2(new_n243), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n256), .B(new_n258), .C1(new_n232), .C2(new_n238), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n248), .B(KEYINPUT94), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT13), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT96), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT96), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n248), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n254), .A2(new_n263), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n265), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n249), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n250), .A2(new_n270), .A3(new_n263), .A4(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT38), .ZN(new_n273));
  XOR2_X1   g072(.A(G64gat), .B(G92gat), .Z(new_n274));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(KEYINPUT37), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  OR2_X1    g093(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n296));
  AOI21_X1  g095(.A(G190gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n295), .A2(new_n302), .A3(new_n296), .ZN(new_n303));
  AND2_X1   g102(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT67), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(G190gat), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n298), .A2(new_n294), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n297), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT23), .B1(new_n284), .B2(new_n285), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  OR2_X1    g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n289), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n300), .A2(KEYINPUT24), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n319), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT25), .B1(new_n315), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT25), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n314), .A2(new_n289), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n324), .B1(new_n317), .B2(new_n318), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n281), .B1(new_n311), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  INV_X1    g133(.A(G190gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n304), .B2(new_n305), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT66), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n337), .A2(new_n294), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(new_n293), .C1(new_n307), .C2(new_n309), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n330), .A2(new_n312), .A3(new_n323), .A4(new_n314), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n340), .A2(KEYINPUT25), .B1(new_n330), .B2(new_n329), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT74), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n334), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT22), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G211gat), .ZN(new_n349));
  INV_X1    g148(.A(G218gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n350), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT22), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(new_n351), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n344), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n311), .B2(new_n332), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n339), .A2(new_n341), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n333), .A2(new_n342), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n370), .A3(new_n357), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n362), .A2(new_n344), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n278), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n280), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n345), .A2(new_n365), .ZN(new_n380));
  INV_X1    g179(.A(new_n358), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n368), .A2(new_n375), .ZN(new_n383));
  INV_X1    g182(.A(new_n371), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n370), .B1(new_n354), .B2(new_n357), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n279), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n273), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n377), .A2(KEYINPUT37), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n278), .B1(new_n366), .B2(new_n376), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(KEYINPUT38), .C1(new_n391), .C2(new_n280), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(G134gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G113gat), .B(G120gat), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n396), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n397));
  INV_X1    g196(.A(G127gat), .ZN(new_n398));
  INV_X1    g197(.A(G120gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G113gat), .ZN(new_n400));
  INV_X1    g199(.A(G113gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G120gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n395), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G141gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(G148gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT79), .B(G141gat), .ZN(new_n410));
  INV_X1    g209(.A(G148gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413));
  OR2_X1    g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(KEYINPUT2), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n411), .A2(G141gat), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n414), .A2(new_n413), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n412), .A2(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(G127gat), .B1(new_n396), .B2(KEYINPUT1), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n398), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(G134gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT4), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n407), .A2(KEYINPUT79), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G141gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n411), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n415), .B1(new_n432), .B2(new_n408), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n406), .A2(new_n423), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n428), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n394), .B(new_n426), .C1(new_n440), .C2(new_n425), .ZN(new_n441));
  INV_X1    g240(.A(new_n420), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT81), .A3(new_n424), .ZN(new_n444));
  INV_X1    g243(.A(new_n394), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n446), .A3(new_n442), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(KEYINPUT5), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n425), .A2(new_n427), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n438), .A2(new_n439), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n424), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT0), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G57gat), .ZN(new_n460));
  INV_X1    g259(.A(G85gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n463), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n462), .A3(new_n456), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n462), .B1(new_n449), .B2(new_n456), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT6), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n465), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n366), .A2(new_n376), .A3(new_n278), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n393), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(G22gat), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n373), .B1(new_n420), .B2(new_n434), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT85), .B1(new_n386), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT29), .B1(new_n354), .B2(new_n357), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n434), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n442), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n372), .B(new_n486), .C1(new_n436), .C2(new_n373), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(G228gat), .A2(G233gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n357), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n355), .B(KEYINPUT83), .C1(new_n356), .C2(new_n351), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n494), .A2(new_n354), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n434), .B1(new_n496), .B2(new_n373), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n497), .B2(new_n442), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n381), .B1(new_n436), .B2(new_n373), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n490), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n492), .B1(new_n490), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n478), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n490), .A2(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n491), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n492), .A3(new_n500), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n477), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n366), .A2(new_n376), .A3(new_n278), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n391), .B1(new_n509), .B2(KEYINPUT30), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n474), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n474), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n454), .A2(new_n445), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n444), .A2(new_n447), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n394), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT39), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n462), .B1(new_n517), .B2(KEYINPUT39), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT40), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n522), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT40), .B1(new_n525), .B2(new_n520), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n524), .A2(new_n526), .A3(new_n470), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n508), .B1(new_n516), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n475), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G71gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G99gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G227gat), .A2(G233gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n421), .A2(new_n422), .A3(G134gat), .ZN(new_n535));
  AOI21_X1  g334(.A(G134gat), .B1(new_n421), .B2(new_n422), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n339), .A2(new_n537), .A3(new_n341), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n339), .B2(new_n341), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n532), .B1(new_n540), .B2(KEYINPUT32), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT69), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n439), .B1(new_n311), .B2(new_n332), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n339), .A2(new_n537), .A3(new_n341), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n533), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n542), .B1(new_n545), .B2(KEYINPUT33), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT33), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(KEYINPUT69), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT70), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n541), .A2(new_n546), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n532), .A2(new_n547), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT34), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n543), .A2(new_n558), .A3(new_n533), .A4(new_n544), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n559), .A2(KEYINPUT71), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n533), .A3(new_n544), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT34), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(KEYINPUT71), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n553), .A2(new_n556), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(KEYINPUT36), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n566), .B1(new_n553), .B2(new_n556), .ZN(new_n570));
  INV_X1    g369(.A(new_n556), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n571), .B(new_n564), .C1(new_n550), .C2(new_n552), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n465), .A2(new_n469), .A3(new_n472), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(new_n510), .A3(new_n513), .A4(new_n515), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n508), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n529), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT86), .ZN(new_n580));
  NOR4_X1   g379(.A1(new_n570), .A2(new_n572), .A3(new_n580), .A4(new_n508), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n473), .A2(new_n516), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n508), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n565), .A2(KEYINPUT86), .A3(new_n584), .A4(new_n567), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n585), .A2(new_n576), .A3(KEYINPUT35), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n578), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  OR2_X1    g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT98), .B(G57gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n593), .A2(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(G57gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(G64gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n589), .B(new_n590), .C1(new_n598), .C2(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n257), .A2(new_n588), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n238), .B1(new_n602), .B2(KEYINPUT21), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n588), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n609), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  OR2_X1    g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G92gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(KEYINPUT8), .A2(new_n618), .B1(new_n461), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n621), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n618), .A3(new_n617), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n623), .A3(new_n622), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n245), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n243), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n630), .B2(new_n602), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n602), .A2(new_n622), .A3(new_n626), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n627), .A2(KEYINPUT103), .A3(new_n600), .A4(new_n624), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G230gat), .ZN(new_n647));
  INV_X1    g446(.A(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n643), .A2(new_n653), .A3(new_n644), .A4(new_n645), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  INV_X1    g457(.A(G176gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n652), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n650), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n614), .A2(new_n641), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT105), .ZN(new_n673));
  AND4_X1   g472(.A1(new_n272), .A2(new_n587), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n473), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g475(.A1(new_n674), .A2(new_n516), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n234), .B2(new_n237), .ZN(new_n678));
  NOR2_X1   g477(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n237), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT42), .B2(new_n680), .ZN(G1325gat));
  NOR2_X1   g482(.A1(new_n570), .A2(new_n572), .ZN(new_n684));
  AOI21_X1  g483(.A(G15gat), .B1(new_n674), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n574), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n685), .B1(new_n674), .B2(new_n687), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n674), .A2(new_n508), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n636), .B(new_n639), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n587), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT35), .B1(new_n585), .B2(new_n576), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n570), .A2(new_n572), .A3(new_n508), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n698), .A2(new_n582), .A3(KEYINPUT86), .A4(new_n579), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n641), .B1(new_n700), .B2(new_n578), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n692), .A3(KEYINPUT44), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n272), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n614), .A3(new_n667), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n575), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n701), .A2(new_n705), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n211), .A3(new_n473), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n212), .A3(new_n516), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT107), .B2(KEYINPUT46), .ZN(new_n713));
  NAND2_X1  g512(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n713), .B(new_n714), .Z(new_n715));
  INV_X1    g514(.A(new_n516), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1329gat));
  NAND2_X1  g517(.A1(new_n686), .A2(G43gat), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n708), .A2(new_n684), .ZN(new_n720));
  OAI22_X1  g519(.A1(new_n706), .A2(new_n719), .B1(G43gat), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g521(.A1(new_n508), .A2(G50gat), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n708), .A2(new_n508), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n706), .A2(new_n723), .B1(G50gat), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g525(.A(new_n272), .B1(new_n700), .B2(new_n578), .ZN(new_n727));
  INV_X1    g526(.A(new_n614), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n693), .A3(new_n668), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n575), .B(KEYINPUT108), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(new_n593), .Z(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(KEYINPUT109), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n727), .A2(KEYINPUT109), .A3(new_n729), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(new_n516), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  AND2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n737), .B2(new_n738), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n730), .A2(new_n684), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(G71gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n686), .B1(new_n734), .B2(new_n735), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G71gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n736), .A2(new_n508), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g548(.A1(new_n614), .A2(new_n272), .A3(new_n668), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n703), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n575), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n614), .A2(new_n272), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n587), .A2(new_n693), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n701), .B2(new_n754), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n461), .A3(new_n473), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n752), .B1(new_n763), .B2(new_n668), .ZN(G1336gat));
  NAND4_X1  g563(.A1(new_n696), .A2(new_n516), .A3(new_n702), .A4(new_n750), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n716), .A2(G92gat), .A3(new_n668), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n759), .B2(new_n761), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n701), .A2(KEYINPUT51), .A3(new_n754), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n765), .A2(G92gat), .B1(new_n773), .B2(new_n769), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n768), .A2(new_n771), .B1(new_n774), .B2(new_n767), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT112), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  OAI221_X1 g576(.A(new_n777), .B1(new_n774), .B2(new_n767), .C1(new_n768), .C2(new_n771), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n751), .B2(new_n574), .ZN(new_n780));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n781), .A3(new_n684), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n668), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n703), .A2(new_n508), .A3(new_n750), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n668), .A2(new_n584), .A3(G106gat), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n762), .A2(new_n788), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n784), .A2(G106gat), .B1(new_n773), .B2(new_n788), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n787), .A2(new_n789), .B1(new_n790), .B2(new_n786), .ZN(G1339gat));
  INV_X1    g590(.A(new_n698), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n663), .B1(new_n656), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n654), .A2(new_n649), .A3(new_n655), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n656), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n664), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n272), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n246), .A2(new_n248), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n259), .A2(new_n261), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n208), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n267), .B2(new_n210), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n668), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n693), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n801), .ZN(new_n809));
  NOR4_X1   g608(.A1(new_n641), .A2(new_n809), .A3(new_n806), .A4(new_n799), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n728), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n672), .A2(new_n704), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n792), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n516), .A2(new_n575), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n704), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n813), .A2(new_n817), .A3(new_n731), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n813), .B2(new_n731), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n716), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n272), .A2(new_n401), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT114), .Z(new_n822));
  OAI21_X1  g621(.A(new_n816), .B1(new_n820), .B2(new_n822), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n815), .B2(new_n668), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n667), .A2(new_n399), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n820), .B2(new_n825), .ZN(G1341gat));
  NOR3_X1   g625(.A1(new_n815), .A2(new_n398), .A3(new_n728), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n820), .A2(new_n728), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n398), .ZN(G1342gat));
  OAI211_X1 g628(.A(new_n693), .B(new_n716), .C1(new_n818), .C2(new_n819), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT56), .B1(new_n830), .B2(G134gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT115), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n830), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n834), .B(KEYINPUT56), .C1(new_n830), .C2(G134gat), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n815), .B2(new_n641), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n574), .A2(new_n814), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n797), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n794), .B(KEYINPUT116), .C1(new_n796), .C2(new_n656), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n798), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n272), .A2(new_n800), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n693), .B1(new_n843), .B2(new_n807), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n728), .B1(new_n844), .B2(new_n810), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n812), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n508), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n838), .B1(new_n847), .B2(KEYINPUT57), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n584), .B1(new_n811), .B2(new_n812), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n272), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n410), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n686), .A2(new_n516), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n731), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(G141gat), .A3(new_n704), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n848), .B2(new_n851), .ZN(new_n860));
  INV_X1    g659(.A(new_n838), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n584), .B1(new_n845), .B2(new_n812), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n850), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT57), .B(new_n584), .C1(new_n811), .C2(new_n812), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n863), .A2(KEYINPUT117), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n272), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n856), .B1(new_n866), .B2(new_n410), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n858), .B1(new_n867), .B2(new_n868), .ZN(G1344gat));
  NOR3_X1   g668(.A1(new_n855), .A2(G148gat), .A3(new_n668), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT118), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT117), .B1(new_n863), .B2(new_n864), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n873), .A2(new_n859), .A3(new_n851), .A4(new_n861), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n411), .C1(new_n875), .C2(new_n667), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n849), .A2(new_n850), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n673), .A2(new_n704), .A3(new_n671), .ZN(new_n879));
  INV_X1    g678(.A(new_n845), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n850), .B(new_n508), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n667), .A3(new_n861), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n871), .B1(new_n876), .B2(new_n884), .ZN(G1345gat));
  INV_X1    g684(.A(new_n855), .ZN(new_n886));
  AOI21_X1  g685(.A(G155gat), .B1(new_n886), .B2(new_n614), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n614), .A2(G155gat), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT119), .Z(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n875), .B2(new_n889), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n886), .B2(new_n693), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n641), .B1(new_n872), .B2(new_n874), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(G162gat), .ZN(G1347gat));
  NAND2_X1  g692(.A1(new_n811), .A2(new_n812), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT120), .B1(new_n894), .B2(new_n575), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n896), .B(new_n473), .C1(new_n811), .C2(new_n812), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n516), .B(new_n698), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(G169gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n272), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n731), .A2(new_n716), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n813), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(new_n272), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n900), .B2(new_n904), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n899), .B2(new_n667), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n668), .A2(new_n659), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n903), .B2(new_n907), .ZN(G1349gat));
  NAND2_X1  g707(.A1(new_n303), .A2(new_n306), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n898), .A2(new_n728), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  INV_X1    g712(.A(new_n903), .ZN(new_n914));
  OAI21_X1  g713(.A(G183gat), .B1(new_n914), .B2(new_n728), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n912), .A2(KEYINPUT121), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT60), .B1(new_n917), .B2(new_n911), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1350gat));
  AOI21_X1  g718(.A(new_n335), .B1(new_n903), .B2(new_n693), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT61), .Z(new_n921));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n335), .A3(new_n693), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1351gat));
  NAND3_X1  g722(.A1(new_n574), .A2(new_n516), .A3(new_n508), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n895), .B2(new_n897), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(G197gat), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n926), .A2(new_n704), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n902), .A2(new_n574), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n882), .A2(new_n272), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n928), .B2(new_n934), .ZN(G1352gat));
  INV_X1    g734(.A(new_n925), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n894), .A2(new_n575), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n896), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n894), .A2(KEYINPUT120), .A3(new_n575), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n661), .A4(new_n667), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n661), .B(new_n925), .C1(new_n895), .C2(new_n897), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT125), .B1(new_n943), .B2(new_n668), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n942), .B2(new_n944), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n882), .A2(new_n667), .A3(new_n932), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n946), .A2(new_n947), .B1(new_n661), .B2(new_n948), .ZN(G1353gat));
  NAND4_X1  g748(.A1(new_n878), .A2(new_n881), .A3(new_n614), .A4(new_n932), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G211gat), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n349), .A3(new_n614), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n951), .A2(new_n957), .A3(new_n952), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n940), .B2(new_n693), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n882), .A2(new_n932), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n641), .A2(new_n350), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1355gat));
endmodule


