//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n464), .B2(KEYINPUT72), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT72), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT71), .B(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n466), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT73), .ZN(G160));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n471), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  INV_X1    g062(.A(new_n473), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n471), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n483), .B1(new_n485), .B2(new_n486), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT74), .Z(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n495), .B1(new_n502), .B2(new_n471), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT3), .B(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n506), .B2(new_n488), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT76), .B(G51), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n522), .A2(G543), .A3(new_n523), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n519), .A2(new_n512), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n532), .A2(G89), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  AND3_X1   g114(.A1(new_n522), .A2(G543), .A3(new_n527), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G52), .B1(G90), .B2(new_n532), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n512), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n515), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n541), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n540), .A2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n532), .A2(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n540), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n512), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n532), .A2(G91), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n540), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n532), .A2(G87), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n512), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n513), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n519), .ZN(G305));
  AOI22_X1  g154(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n515), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n532), .A2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n540), .A2(G47), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(new_n581), .B2(new_n582), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n585), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n532), .A2(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n522), .A2(G543), .A3(new_n527), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n592), .A2(new_n515), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G321));
  AND2_X1   g176(.A1(new_n562), .A2(new_n566), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT81), .B1(new_n602), .B2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  MUX2_X1   g179(.A(KEYINPUT81), .B(new_n603), .S(new_n604), .Z(G297));
  MUX2_X1   g180(.A(KEYINPUT81), .B(new_n603), .S(new_n604), .Z(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n599), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g186(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n612));
  XNOR2_X1  g187(.A(G323), .B(new_n612), .ZN(G282));
  NAND2_X1  g188(.A1(new_n505), .A2(new_n465), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  INV_X1    g192(.A(new_n485), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G135), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n489), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n473), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n622), .A2(G123), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n617), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT86), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n638), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  MUX2_X1   g246(.A(new_n671), .B(new_n670), .S(new_n663), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G25), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n622), .A2(G119), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n618), .A2(G131), .ZN(new_n684));
  OAI221_X1 g259(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n473), .C2(G107), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n686), .B2(G29), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT88), .Z(new_n690));
  XOR2_X1   g265(.A(KEYINPUT89), .B(G16), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G24), .B(G290), .S(new_n692), .Z(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G1986), .Z(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT92), .Z(new_n702));
  MUX2_X1   g277(.A(G6), .B(G305), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT32), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1981), .Z(new_n705));
  NOR2_X1   g280(.A1(new_n692), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n692), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1971), .Z(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n690), .B(new_n694), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n710), .B2(new_n709), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT36), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n555), .A2(new_n692), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G19), .B2(new_n692), .ZN(new_n715));
  INV_X1    g290(.A(G1341), .ZN(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  NAND2_X1  g292(.A1(G164), .A2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G27), .B2(G29), .ZN(new_n719));
  OAI22_X1  g294(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT25), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n505), .A2(G127), .ZN(new_n726));
  INV_X1    g301(.A(G115), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n464), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n488), .A2(new_n728), .B1(new_n618), .B2(G139), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n724), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G33), .B(new_n730), .S(G29), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2072), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n720), .B(new_n732), .C1(new_n717), .C2(new_n719), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n627), .A2(new_n680), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT26), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n737), .A2(new_n738), .B1(G105), .B2(new_n465), .ZN(new_n739));
  INV_X1    g314(.A(G141), .ZN(new_n740));
  INV_X1    g315(.A(G129), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n739), .B1(new_n485), .B2(new_n740), .C1(new_n489), .C2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G32), .B(new_n742), .S(G29), .Z(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G11), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G28), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n680), .B1(new_n749), .B2(G28), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n747), .B(new_n748), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n734), .A2(new_n745), .A3(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n715), .A2(new_n716), .B1(new_n743), .B2(new_n744), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n695), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n695), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G1961), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n680), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  OAI221_X1 g334(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  INV_X1    g336(.A(G128), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n760), .B1(new_n485), .B2(new_n761), .C1(new_n762), .C2(new_n489), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n759), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2067), .ZN(new_n765));
  AND4_X1   g340(.A1(new_n753), .A2(new_n754), .A3(new_n757), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n680), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n680), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n733), .B(new_n766), .C1(G2090), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(G160), .A2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n773), .B2(KEYINPUT24), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(KEYINPUT24), .B2(new_n773), .ZN(new_n775));
  AOI21_X1  g350(.A(G2084), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n772), .A2(G2084), .A3(new_n775), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n776), .B(new_n777), .C1(G1961), .C2(new_n756), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n695), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n695), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n691), .A2(G20), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT95), .B(KEYINPUT23), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1956), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n780), .A2(G1966), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n778), .A2(new_n781), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n770), .A2(G2090), .ZN(new_n789));
  NOR2_X1   g364(.A1(G4), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n599), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1348), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n771), .A2(new_n788), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n713), .A2(new_n793), .ZN(G150));
  INV_X1    g369(.A(G150), .ZN(G311));
  NAND2_X1  g370(.A1(new_n532), .A2(G93), .ZN(new_n796));
  INV_X1    g371(.A(G55), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n796), .B1(new_n593), .B2(new_n797), .C1(new_n798), .C2(new_n515), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G860), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT37), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n599), .A2(G559), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT38), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n554), .B(new_n799), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT97), .ZN(new_n808));
  INV_X1    g383(.A(G860), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n806), .B2(KEYINPUT39), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n801), .B1(new_n808), .B2(new_n810), .ZN(G145));
  AOI22_X1  g386(.A1(new_n622), .A2(G130), .B1(new_n618), .B2(G142), .ZN(new_n812));
  INV_X1    g387(.A(G118), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n488), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(new_n615), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n686), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT99), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n763), .B(new_n508), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n730), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n742), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n627), .B(G160), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n491), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(G37), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(KEYINPUT100), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n824), .A2(new_n820), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n830), .B(new_n831), .C1(new_n824), .C2(new_n821), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n835));
  INV_X1    g410(.A(new_n599), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(new_n602), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n599), .A2(G299), .A3(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n602), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(KEYINPUT102), .A3(new_n838), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n609), .B(new_n805), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n841), .A2(KEYINPUT41), .A3(new_n842), .A4(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n839), .A2(new_n842), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT41), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n845), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(G290), .B(G305), .Z(new_n854));
  XNOR2_X1  g429(.A(G166), .B(G288), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n854), .B(new_n855), .Z(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT42), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n853), .B(new_n857), .ZN(new_n858));
  MUX2_X1   g433(.A(new_n799), .B(new_n858), .S(G868), .Z(G295));
  MUX2_X1   g434(.A(new_n799), .B(new_n858), .S(G868), .Z(G331));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n848), .A2(new_n851), .ZN(new_n862));
  OAI21_X1  g437(.A(G168), .B1(G301), .B2(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g438(.A1(G301), .A2(KEYINPUT104), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n863), .B(new_n864), .Z(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(new_n805), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n805), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n839), .A2(new_n840), .B1(new_n602), .B2(new_n836), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n870), .B2(new_n843), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n865), .A2(KEYINPUT105), .A3(new_n805), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT105), .B1(new_n865), .B2(new_n805), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n862), .A2(new_n869), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n856), .ZN(new_n876));
  OAI211_X1 g451(.A(KEYINPUT106), .B(new_n861), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n862), .A2(new_n869), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n874), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n871), .A2(new_n874), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n848), .A2(new_n851), .B1(new_n868), .B2(new_n867), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n856), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT106), .B1(new_n884), .B2(new_n861), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n875), .B2(new_n876), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n841), .A2(new_n850), .A3(new_n842), .A4(new_n843), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n849), .A2(KEYINPUT41), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n872), .A2(new_n873), .A3(new_n866), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n844), .A2(new_n867), .ZN(new_n893));
  INV_X1    g468(.A(new_n868), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n891), .A2(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n856), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n887), .A2(KEYINPUT107), .A3(new_n888), .A4(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n888), .A3(new_n861), .A4(new_n880), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n886), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n888), .B1(new_n881), .B2(new_n885), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n887), .A2(KEYINPUT43), .A3(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n901), .B(new_n904), .S(KEYINPUT44), .Z(G397));
  INV_X1    g480(.A(G1384), .ZN(new_n906));
  INV_X1    g481(.A(new_n495), .ZN(new_n907));
  INV_X1    g482(.A(new_n501), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n473), .B2(new_n499), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n909), .B2(new_n472), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n476), .A2(new_n477), .A3(G138), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT4), .B1(new_n911), .B2(new_n473), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n906), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n496), .A2(new_n498), .A3(G137), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n916), .A2(new_n471), .B1(G101), .B2(new_n465), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n478), .A2(new_n479), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n917), .B(G40), .C1(new_n918), .C2(new_n473), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n921), .A2(G290), .A3(G1986), .ZN(new_n922));
  AND3_X1   g497(.A1(G290), .A2(G1986), .A3(new_n920), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(G2067), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n763), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n742), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n686), .B(new_n688), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n921), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT117), .ZN(new_n935));
  XNOR2_X1  g510(.A(G299), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT116), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT57), .B1(new_n562), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n936), .B(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n919), .B1(new_n913), .B2(KEYINPUT50), .ZN(new_n940));
  NOR2_X1   g515(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n910), .B2(new_n912), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT115), .B(G1956), .Z(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n503), .B2(new_n507), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n475), .A2(new_n948), .A3(new_n480), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n915), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT56), .B(G2072), .Z(new_n951));
  OAI21_X1  g526(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n939), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n949), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n942), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n508), .A2(KEYINPUT109), .A3(new_n941), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1348), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n949), .A2(new_n946), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n960), .A2(new_n961), .B1(new_n926), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(new_n836), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n953), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n939), .A2(new_n952), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n953), .A2(new_n967), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT60), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n972), .A3(new_n599), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n967), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n964), .A2(new_n836), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT60), .B1(new_n975), .B2(new_n965), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n971), .A2(new_n973), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT58), .B(G1341), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n950), .A2(G1996), .B1(new_n963), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n555), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  NOR2_X1   g557(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n982), .B(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n968), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(G305), .B(G1981), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT49), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n962), .A2(G8), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(G288), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n697), .B2(G1976), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n992), .A2(KEYINPUT52), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n950), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G1971), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT110), .B(G2090), .Z(new_n1002));
  NOR2_X1   g577(.A1(new_n943), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G8), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n960), .A2(new_n1002), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1008), .B2(new_n1001), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(new_n1006), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n999), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n950), .A2(G2078), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(KEYINPUT53), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(KEYINPUT53), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n959), .A2(G1961), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(G301), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(G301), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1012), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT109), .B1(new_n508), .B2(new_n941), .ZN(new_n1025));
  INV_X1    g600(.A(new_n941), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n956), .B(new_n1026), .C1(new_n503), .C2(new_n507), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n940), .B(new_n1024), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n950), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n957), .A2(new_n958), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(KEYINPUT113), .A3(new_n1024), .A4(new_n940), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n537), .B2(new_n538), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT120), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(G8), .C1(new_n537), .C2(new_n538), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT113), .B1(new_n959), .B2(new_n1024), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1034), .A2(new_n1032), .ZN(new_n1043));
  OAI21_X1  g618(.A(G8), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1039), .A4(new_n1037), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1037), .A2(KEYINPUT122), .A3(new_n1039), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT122), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1035), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1046), .B1(new_n1053), .B2(KEYINPUT123), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1055), .B(new_n1045), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1041), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT124), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1041), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1023), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n986), .B1(new_n1061), .B2(KEYINPUT125), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1063), .B(new_n1023), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1060), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1035), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT121), .B1(new_n1035), .B2(G8), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1049), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1055), .B1(new_n1069), .B2(new_n1045), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1053), .A2(KEYINPUT123), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1046), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1059), .B1(new_n1072), .B2(new_n1041), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1058), .A2(new_n1075), .A3(new_n1060), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(G1976), .B(G288), .C1(new_n988), .C2(new_n989), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G305), .A2(G1981), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n989), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n999), .B(KEYINPUT112), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1010), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1009), .A2(new_n1006), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1010), .A2(KEYINPUT63), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1044), .A2(G286), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1087), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1011), .B2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1086), .A2(new_n1087), .B1(KEYINPUT114), .B2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1090), .A2(KEYINPUT114), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1083), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1078), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n934), .B1(new_n1065), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n922), .A2(KEYINPUT48), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n922), .A2(KEYINPUT48), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n933), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n920), .A2(new_n928), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT46), .ZN(new_n1100));
  INV_X1    g675(.A(new_n927), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n920), .B1(new_n1101), .B2(new_n742), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT47), .Z(new_n1104));
  NAND4_X1  g679(.A1(new_n683), .A2(new_n684), .A3(new_n688), .A4(new_n685), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n930), .A2(new_n1105), .B1(G2067), .B2(new_n763), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1098), .B(new_n1104), .C1(new_n920), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1095), .A2(new_n1107), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g683(.A1(G227), .A2(new_n462), .ZN(new_n1110));
  NAND2_X1  g684(.A1(new_n648), .A2(new_n1110), .ZN(new_n1111));
  OR3_X1    g685(.A1(G229), .A2(new_n1111), .A3(KEYINPUT126), .ZN(new_n1112));
  OAI21_X1  g686(.A(KEYINPUT126), .B1(G229), .B2(new_n1111), .ZN(new_n1113));
  AOI22_X1  g687(.A1(new_n1112), .A2(new_n1113), .B1(new_n829), .B2(new_n832), .ZN(new_n1114));
  INV_X1    g688(.A(KEYINPUT127), .ZN(new_n1115));
  AND2_X1   g689(.A1(new_n877), .A2(new_n880), .ZN(new_n1116));
  NAND2_X1  g690(.A1(new_n884), .A2(new_n861), .ZN(new_n1117));
  INV_X1    g691(.A(KEYINPUT106), .ZN(new_n1118));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g693(.A(new_n888), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g694(.A1(new_n900), .A2(new_n897), .ZN(new_n1121));
  OAI211_X1 g695(.A(new_n1114), .B(new_n1115), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g696(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n901), .B2(new_n1114), .ZN(new_n1124));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n1124), .ZN(G308));
  NAND2_X1  g699(.A1(new_n901), .A2(new_n1114), .ZN(G225));
endmodule


