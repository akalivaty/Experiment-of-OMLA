//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT68), .ZN(new_n204));
  XOR2_X1   g003(.A(G71gat), .B(G99gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(G127gat), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n208), .A2(KEYINPUT1), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(G113gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G120gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n223), .B(new_n224), .C1(new_n227), .C2(new_n222), .ZN(new_n228));
  OR2_X1    g027(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT27), .B(G183gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n231), .A2(KEYINPUT67), .A3(KEYINPUT28), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n234), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  OR3_X1    g041(.A1(new_n238), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT27), .B1(new_n238), .B2(KEYINPUT66), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n231), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n228), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n225), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n229), .A2(new_n230), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(G183gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n252), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n258), .A2(new_n259), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n221), .B1(new_n248), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n262), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n259), .B1(new_n252), .B2(new_n257), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n212), .A2(new_n220), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n241), .A2(new_n233), .B1(new_n245), .B2(new_n246), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n269), .B(new_n270), .C1(new_n271), .C2(new_n228), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n207), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n266), .A2(new_n272), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT34), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT34), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n266), .A2(new_n272), .A3(new_n281), .A4(new_n274), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n274), .B1(new_n266), .B2(new_n272), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n206), .B1(new_n287), .B2(KEYINPUT33), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n280), .A3(new_n282), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n284), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n202), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n285), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT36), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G211gat), .B(G218gat), .Z(new_n298));
  AOI21_X1  g097(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n299));
  AND2_X1   g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n305), .C1(new_n301), .C2(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT69), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n298), .B(new_n309), .C1(new_n299), .C2(new_n302), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314));
  OR2_X1    g113(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n321), .ZN(new_n327));
  NAND2_X1  g126(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n329), .B2(G162gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G155gat), .B(G162gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n314), .A3(new_n316), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n324), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G228gat), .ZN(new_n335));
  INV_X1    g134(.A(G233gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n307), .A2(new_n338), .A3(new_n310), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n307), .B2(new_n310), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n324), .B(new_n312), .C1(new_n330), .C2(new_n332), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n347));
  OAI21_X1  g146(.A(G162gat), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT2), .ZN(new_n349));
  AND4_X1   g148(.A1(new_n320), .A2(new_n314), .A3(new_n322), .A4(new_n316), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n349), .A2(new_n350), .B1(new_n323), .B2(new_n318), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT74), .A3(new_n312), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n334), .B(new_n337), .C1(new_n342), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n303), .A2(new_n306), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n308), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n356), .B2(new_n312), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n308), .ZN(new_n359));
  INV_X1    g158(.A(new_n341), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n339), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n362), .B2(new_n337), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G22gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT31), .B(G50gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G22gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n354), .B(new_n369), .C1(new_n362), .C2(new_n337), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n364), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  INV_X1    g171(.A(new_n357), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n342), .B2(new_n353), .ZN(new_n374));
  INV_X1    g173(.A(new_n337), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n361), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n313), .B2(new_n333), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n374), .A2(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n378), .B2(new_n369), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT81), .A3(G22gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n375), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n383), .A2(KEYINPUT80), .A3(new_n369), .A4(new_n354), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n379), .A2(new_n380), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n371), .B1(new_n385), .B2(new_n367), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT0), .ZN(new_n388));
  XNOR2_X1  g187(.A(G57gat), .B(G85gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  NOR2_X1   g189(.A1(new_n333), .A2(new_n221), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n333), .B2(new_n221), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n270), .A2(new_n351), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(KEYINPUT4), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n270), .B1(new_n333), .B2(KEYINPUT3), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT75), .B1(new_n358), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n402), .B(KEYINPUT76), .Z(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n390), .B1(new_n404), .B2(KEYINPUT39), .ZN(new_n405));
  INV_X1    g204(.A(new_n403), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT74), .B1(new_n351), .B2(new_n312), .ZN(new_n407));
  XOR2_X1   g206(.A(G141gat), .B(G148gat), .Z(new_n408));
  AOI21_X1  g207(.A(new_n319), .B1(new_n327), .B2(new_n328), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n331), .B(new_n408), .C1(new_n409), .C2(new_n325), .ZN(new_n410));
  AND4_X1   g209(.A1(KEYINPUT74), .A2(new_n410), .A3(new_n312), .A4(new_n324), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n398), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT75), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n398), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n406), .B1(new_n416), .B2(new_n397), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n393), .B(new_n395), .C1(new_n351), .C2(new_n270), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n418), .A2(new_n403), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT39), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n403), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n397), .B(new_n425), .C1(new_n399), .C2(new_n400), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n395), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n403), .B1(new_n391), .B2(KEYINPUT4), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n414), .B2(new_n415), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n418), .A2(new_n403), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n424), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n428), .A2(new_n429), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n399), .B2(new_n400), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n423), .B1(new_n418), .B2(new_n403), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT79), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n426), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n390), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n422), .A2(KEYINPUT40), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT71), .ZN(new_n444));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n269), .B1(new_n271), .B2(new_n228), .ZN(new_n448));
  NAND2_X1  g247(.A1(G226gat), .A2(G233gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n448), .B2(new_n308), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(new_n342), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n248), .A2(new_n265), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n455), .B2(KEYINPUT29), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n361), .B1(new_n456), .B2(new_n451), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n447), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n342), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n361), .A3(new_n451), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n446), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n447), .C1(new_n454), .C2(new_n457), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n441), .B1(new_n417), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n404), .A2(KEYINPUT39), .A3(new_n419), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT40), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n386), .B1(new_n442), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n440), .A2(new_n441), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n390), .B(new_n426), .C1(new_n435), .C2(new_n439), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n426), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n434), .B1(new_n431), .B2(new_n433), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n437), .A2(KEYINPUT79), .A3(new_n438), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n479), .A2(new_n473), .A3(new_n390), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n460), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(new_n459), .B2(new_n460), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT38), .B(new_n446), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n485), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n447), .B1(new_n487), .B2(new_n483), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n458), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n481), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n297), .B1(new_n471), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n473), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n390), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n465), .B1(new_n496), .B2(new_n480), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n386), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n290), .A2(new_n291), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n385), .A2(new_n367), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n502), .B(new_n503), .C1(new_n504), .C2(new_n371), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n501), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n294), .A2(new_n295), .ZN(new_n507));
  INV_X1    g306(.A(new_n503), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n386), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n475), .A2(new_n481), .ZN(new_n510));
  INV_X1    g309(.A(new_n501), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n509), .A2(new_n510), .A3(new_n465), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n499), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  INV_X1    g314(.A(G15gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(G22gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n369), .A2(G15gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n369), .A2(G15gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(G22gat), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT16), .B1(KEYINPUT83), .B2(G1gat), .ZN(new_n522));
  AND2_X1   g321(.A1(KEYINPUT83), .A2(G1gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n522), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n521), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n529), .A3(G8gat), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n519), .B(new_n524), .C1(new_n526), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  AND2_X1   g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(KEYINPUT14), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G43gat), .B(G50gat), .Z(new_n538));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT15), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT15), .B1(new_n537), .B2(new_n540), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT14), .ZN(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n540), .A3(KEYINPUT15), .A4(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G43gat), .B(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n534), .B(new_n541), .C1(new_n542), .C2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n540), .A3(new_n546), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n547), .A3(new_n548), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n534), .B1(new_n555), .B2(new_n541), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n533), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n530), .A2(new_n532), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n541), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT85), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n561), .A2(new_n562), .B1(G229gat), .B2(G233gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n557), .A2(new_n560), .A3(new_n567), .A4(new_n563), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n530), .A2(new_n555), .A3(new_n532), .A4(new_n541), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n547), .A2(new_n548), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n547), .A2(new_n548), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n554), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT87), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n532), .A4(new_n530), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n560), .A2(KEYINPUT86), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT86), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n558), .A2(new_n579), .A3(new_n559), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT13), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G197gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT11), .B(G169gat), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n589), .A2(KEYINPUT12), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT12), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n581), .B2(new_n583), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT88), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n569), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n569), .B2(new_n595), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n514), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n603), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n603), .A3(new_n609), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT95), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n605), .A2(new_n603), .A3(new_n609), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n556), .B2(new_n551), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n602), .A2(KEYINPUT97), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n617), .B2(new_n574), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI211_X1 g423(.A(KEYINPUT97), .B(new_n602), .C1(new_n620), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n624), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n602), .A2(KEYINPUT97), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n625), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n625), .B2(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  INV_X1    g435(.A(G71gat), .ZN(new_n637));
  INV_X1    g436(.A(G78gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT9), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT91), .B(G57gat), .ZN(new_n642));
  INV_X1    g441(.A(G64gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(G57gat), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(G71gat), .A2(G78gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(G71gat), .A2(G78gat), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT89), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT89), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n639), .A2(new_n650), .A3(new_n636), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT90), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n640), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n643), .A2(G57gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n645), .B2(new_n655), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n652), .B2(new_n656), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n646), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT21), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n533), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT94), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G127gat), .B(G155gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NAND2_X1  g467(.A1(G231gat), .A2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT92), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G183gat), .B(G211gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n666), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n635), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(G230gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n336), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n605), .A2(new_n609), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT98), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n646), .B(new_n680), .C1(new_n657), .C2(new_n658), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n615), .A2(new_n610), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT89), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n650), .B1(new_n639), .B2(new_n636), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n656), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n690), .A2(new_n646), .A3(new_n682), .A4(new_n680), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT10), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT10), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n617), .A2(new_n693), .A3(new_n659), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n678), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n684), .A2(new_n691), .A3(new_n677), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n696), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n696), .B2(new_n698), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n675), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n601), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n510), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(new_n515), .ZN(G1324gat));
  INV_X1    g509(.A(new_n708), .ZN(new_n711));
  INV_X1    g510(.A(new_n465), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n531), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G8gat), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n708), .A2(new_n465), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT42), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT42), .B2(new_n716), .ZN(G1325gat));
  INV_X1    g517(.A(new_n297), .ZN(new_n719));
  OAI21_X1  g518(.A(G15gat), .B1(new_n708), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n502), .A2(new_n516), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n708), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT100), .Z(G1326gat));
  INV_X1    g522(.A(new_n386), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT43), .B(G22gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  NOR2_X1   g526(.A1(new_n674), .A2(new_n706), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n635), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n601), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n510), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n543), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT45), .ZN(new_n734));
  INV_X1    g533(.A(new_n635), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n499), .B2(new_n513), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(KEYINPUT44), .B(new_n735), .C1(new_n499), .C2(new_n513), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n599), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n594), .B(KEYINPUT101), .C1(new_n597), .C2(new_n598), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n740), .A2(new_n510), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n734), .B1(new_n543), .B2(new_n747), .ZN(G1328gat));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n544), .A3(new_n712), .ZN(new_n749));
  AND2_X1   g548(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n740), .A2(new_n465), .A3(new_n746), .ZN(new_n753));
  OAI221_X1 g552(.A(new_n752), .B1(new_n544), .B2(new_n753), .C1(new_n750), .C2(new_n749), .ZN(G1329gat));
  NOR2_X1   g553(.A1(new_n507), .A2(G43gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n731), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n297), .A3(new_n739), .A4(new_n745), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n758), .A3(KEYINPUT47), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n758), .A2(KEYINPUT103), .B1(new_n731), .B2(new_n755), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n761), .A3(G43gat), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT104), .B(KEYINPUT47), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n758), .A2(KEYINPUT103), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n762), .A3(new_n756), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n759), .B1(new_n763), .B2(new_n768), .ZN(G1330gat));
  NAND4_X1  g568(.A1(new_n738), .A2(new_n386), .A3(new_n739), .A4(new_n745), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n770), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n724), .A2(G50gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n601), .A2(new_n730), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n601), .A2(KEYINPUT106), .A3(new_n730), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n770), .A2(G50gat), .B1(KEYINPUT105), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n771), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n773), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT107), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n773), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT48), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n777), .A2(new_n779), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n771), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(G1331gat));
  NAND2_X1  g587(.A1(new_n744), .A2(new_n706), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n514), .A2(new_n675), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n732), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(new_n642), .ZN(G1332gat));
  XNOR2_X1  g591(.A(new_n465), .B(KEYINPUT108), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT109), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1333gat));
  INV_X1    g598(.A(new_n790), .ZN(new_n800));
  OAI21_X1  g599(.A(G71gat), .B1(new_n800), .B2(new_n719), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n790), .A2(new_n637), .A3(new_n502), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n803), .B(new_n804), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n386), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  INV_X1    g606(.A(new_n674), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n744), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n736), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n732), .A2(new_n607), .A3(new_n706), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n789), .A2(new_n674), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n740), .A2(new_n510), .A3(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n814), .A2(new_n815), .B1(new_n607), .B2(new_n818), .ZN(G1336gat));
  NOR3_X1   g618(.A1(new_n740), .A2(new_n794), .A3(new_n817), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(G92gat), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n793), .A2(new_n608), .A3(new_n706), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT111), .Z(new_n827));
  NAND2_X1  g626(.A1(new_n813), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n740), .A2(new_n465), .A3(new_n817), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n608), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1337gat));
  INV_X1    g632(.A(G99gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n502), .A2(new_n834), .A3(new_n706), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n740), .A2(new_n719), .A3(new_n817), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n814), .A2(new_n835), .B1(new_n834), .B2(new_n836), .ZN(G1338gat));
  INV_X1    g636(.A(new_n706), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n724), .A2(G106gat), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n738), .A2(new_n386), .A3(new_n739), .A4(new_n816), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n813), .A2(new_n839), .B1(G106gat), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT113), .B1(new_n840), .B2(G106gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n841), .B(new_n843), .ZN(G1339gat));
  NAND2_X1  g643(.A1(new_n707), .A2(new_n744), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n684), .A2(new_n691), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n693), .ZN(new_n849));
  INV_X1    g648(.A(new_n694), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n847), .B1(new_n851), .B2(new_n678), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n850), .A3(new_n677), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n847), .B(new_n678), .C1(new_n692), .C2(new_n694), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n702), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n846), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n852), .B2(new_n853), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n703), .B1(new_n858), .B2(KEYINPUT55), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n597), .A2(new_n598), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n581), .A2(new_n583), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n582), .B1(new_n557), .B2(new_n560), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n590), .B(new_n589), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n635), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n742), .A2(new_n743), .A3(new_n857), .A4(new_n859), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n706), .A2(new_n861), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n735), .B1(new_n869), .B2(KEYINPUT114), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n866), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n845), .B1(new_n873), .B2(new_n674), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n724), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n732), .A3(new_n502), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n793), .ZN(new_n877));
  INV_X1    g676(.A(new_n744), .ZN(new_n878));
  AOI21_X1  g677(.A(G113gat), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n600), .A2(new_n215), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n877), .B2(new_n880), .ZN(G1340gat));
  NAND2_X1  g680(.A1(KEYINPUT115), .A2(G120gat), .ZN(new_n882));
  XNOR2_X1  g681(.A(KEYINPUT115), .B(G120gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n877), .A2(new_n706), .ZN(new_n884));
  MUX2_X1   g683(.A(new_n882), .B(new_n883), .S(new_n884), .Z(G1341gat));
  NAND2_X1  g684(.A1(new_n877), .A2(new_n674), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g686(.A1(new_n735), .A2(new_n465), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n876), .A2(G134gat), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n876), .A2(new_n635), .A3(new_n793), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n209), .B2(new_n892), .ZN(G1343gat));
  XNOR2_X1  g692(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n635), .A3(new_n872), .ZN(new_n896));
  INV_X1    g695(.A(new_n866), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n674), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n845), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n386), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n297), .A2(new_n510), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n793), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n600), .A2(G141gat), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT118), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n894), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n874), .B2(new_n386), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n724), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n868), .B1(new_n860), .B2(new_n600), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n635), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n808), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n918), .B2(new_n845), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n904), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n910), .B1(new_n920), .B2(new_n600), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G141gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n920), .A2(new_n910), .A3(new_n600), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n909), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n900), .B2(new_n912), .ZN(new_n925));
  INV_X1    g724(.A(new_n904), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT117), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(new_n904), .C1(new_n911), .C2(new_n919), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n878), .A3(new_n929), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n930), .A2(G141gat), .B1(new_n906), .B2(new_n908), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(G1344gat));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n934), .B(G148gat), .C1(new_n906), .C2(new_n706), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n927), .A2(new_n706), .A3(new_n929), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n934), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n874), .A2(new_n913), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n917), .A2(new_n808), .B1(new_n600), .B2(new_n707), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n912), .B1(new_n939), .B2(new_n724), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI211_X1 g740(.A(new_n934), .B(new_n838), .C1(new_n926), .C2(KEYINPUT121), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n941), .B(new_n942), .C1(KEYINPUT121), .C2(new_n926), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n935), .B1(new_n944), .B2(G148gat), .ZN(G1345gat));
  NAND2_X1  g744(.A1(new_n927), .A2(new_n929), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n329), .B1(new_n946), .B2(new_n808), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n674), .A2(new_n327), .A3(new_n328), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n905), .B2(new_n948), .ZN(G1346gat));
  OR4_X1    g748(.A1(G162gat), .A2(new_n900), .A3(new_n888), .A4(new_n903), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT122), .ZN(new_n951));
  OAI21_X1  g750(.A(G162gat), .B1(new_n946), .B2(new_n635), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1347gat));
  NOR3_X1   g752(.A1(new_n732), .A2(new_n465), .A3(new_n507), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n875), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(G169gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(new_n600), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n874), .A2(new_n510), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n794), .A2(new_n386), .A3(new_n507), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n878), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n957), .B1(new_n956), .B2(new_n962), .ZN(G1348gat));
  OAI21_X1  g762(.A(G176gat), .B1(new_n955), .B2(new_n838), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n838), .A2(G176gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n960), .B2(new_n965), .ZN(G1349gat));
  OAI21_X1  g765(.A(G183gat), .B1(new_n955), .B2(new_n808), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n808), .A2(new_n240), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  NOR4_X1   g769(.A1(new_n960), .A2(KEYINPUT123), .A3(new_n240), .A4(new_n808), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT60), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT60), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n974), .B(new_n967), .C1(new_n970), .C2(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n231), .A3(new_n735), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n955), .B2(new_n635), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  NAND3_X1  g780(.A1(new_n719), .A2(new_n386), .A3(new_n793), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT124), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n958), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(G197gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n985), .A2(new_n986), .A3(new_n878), .ZN(new_n987));
  INV_X1    g786(.A(new_n941), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n719), .A2(new_n510), .A3(new_n712), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n988), .A2(new_n600), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n990), .B2(new_n986), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT125), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n987), .B(new_n993), .C1(new_n990), .C2(new_n986), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1352gat));
  XOR2_X1   g794(.A(KEYINPUT126), .B(G204gat), .Z(new_n996));
  NAND3_X1  g795(.A1(new_n985), .A2(new_n706), .A3(new_n996), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n988), .A2(new_n838), .A3(new_n989), .ZN(new_n1000));
  OAI211_X1 g799(.A(new_n998), .B(new_n999), .C1(new_n1000), .C2(new_n996), .ZN(G1353gat));
  OR3_X1    g800(.A1(new_n984), .A2(G211gat), .A3(new_n808), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n988), .A2(new_n989), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(new_n674), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  AOI21_X1  g806(.A(G218gat), .B1(new_n985), .B2(new_n735), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n735), .A2(G218gat), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT127), .Z(new_n1010));
  AOI21_X1  g809(.A(new_n1008), .B1(new_n1003), .B2(new_n1010), .ZN(G1355gat));
endmodule


