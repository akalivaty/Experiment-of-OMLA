//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND2_X1  g026(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n469), .A2(new_n474), .A3(new_n476), .A4(new_n470), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n466), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XOR2_X1   g059(.A(KEYINPUT69), .B(G2105), .Z(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n485), .C2(G112), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n471), .A2(new_n465), .A3(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n474), .A2(new_n476), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n477), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n485), .A2(new_n498), .A3(G138), .A4(new_n465), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  AOI211_X1 g077(.A(new_n502), .B(new_n495), .C1(new_n497), .C2(new_n499), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(G62), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n508), .A2(new_n509), .B1(G75), .B2(G543), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT71), .B(G62), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G50), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n506), .A2(new_n507), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n512), .A2(new_n520), .ZN(G166));
  AOI22_X1  g096(.A1(new_n519), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n514), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(new_n524), .A3(new_n518), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT72), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n525), .A2(new_n528), .A3(G543), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT73), .B(G51), .Z(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n523), .A2(new_n531), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n536));
  INV_X1    g111(.A(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT5), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n519), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n514), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(G90), .A2(new_n541), .B1(new_n544), .B2(G651), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G52), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n529), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n540), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n505), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n529), .A2(G43), .B1(G81), .B2(new_n541), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n514), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(KEYINPUT76), .A3(G651), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(new_n569), .B1(G91), .B2(new_n541), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n525), .A2(new_n528), .A3(G543), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n571), .A2(KEYINPUT9), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n571), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(new_n512), .B2(new_n520), .ZN(new_n578));
  NAND2_X1  g153(.A1(G75), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G62), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n538), .B2(new_n539), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n581), .B2(KEYINPUT71), .ZN(new_n582));
  INV_X1    g157(.A(new_n511), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n516), .A2(new_n519), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(KEYINPUT77), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n578), .A2(new_n586), .ZN(G303));
  NAND4_X1  g162(.A1(new_n525), .A2(new_n528), .A3(G49), .A4(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n519), .A2(new_n540), .A3(G87), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  OAI21_X1  g166(.A(G61), .B1(new_n506), .B2(new_n507), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  OAI21_X1  g170(.A(G86), .B1(new_n506), .B2(new_n507), .ZN(new_n596));
  NAND2_X1  g171(.A1(G48), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n519), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n541), .A2(G85), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT78), .B(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n540), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI221_X1 g178(.A(new_n601), .B1(new_n571), .B2(new_n602), .C1(new_n505), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(KEYINPUT79), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n605), .A2(KEYINPUT79), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n540), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n505), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G54), .B2(new_n529), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n519), .A2(new_n540), .A3(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n606), .B1(new_n607), .B2(new_n615), .ZN(G284));
  AOI21_X1  g191(.A(new_n606), .B1(new_n607), .B2(new_n615), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT80), .Z(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G280));
  INV_X1    g197(.A(new_n613), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT81), .B(G559), .Z(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(G860), .B2(new_n624), .ZN(G148));
  NAND2_X1  g200(.A1(new_n555), .A2(new_n614), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n623), .A2(new_n624), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n483), .A2(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n483), .A2(G135), .ZN(new_n637));
  OAI221_X1 g212(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n485), .C2(G111), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n471), .A2(new_n465), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n644), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(KEYINPUT83), .B1(new_n656), .B2(new_n644), .ZN(new_n660));
  OAI221_X1 g235(.A(G14), .B1(new_n644), .B2(new_n656), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  INV_X1    g245(.A(new_n663), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n666), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT85), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n683), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(KEYINPUT20), .A3(new_n683), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n685), .B1(new_n683), .B2(new_n681), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT86), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n695), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n677), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(new_n676), .A3(new_n696), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G23), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT33), .ZN(new_n708));
  INV_X1    g283(.A(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G22), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G166), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1971), .ZN(new_n713));
  NOR2_X1   g288(.A1(G6), .A2(G16), .ZN(new_n714));
  AOI22_X1  g289(.A1(G651), .A2(new_n594), .B1(new_n598), .B2(new_n519), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT32), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1981), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n710), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1986), .Z(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G25), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n471), .A2(new_n465), .A3(G119), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT87), .Z(new_n728));
  OR2_X1    g303(.A1(new_n485), .A2(G107), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n729), .A2(new_n731), .B1(new_n483), .B2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n726), .B1(new_n734), .B2(new_n725), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n721), .A2(new_n722), .A3(new_n724), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(G19), .ZN(new_n740));
  OR3_X1    g315(.A1(new_n740), .A2(KEYINPUT88), .A3(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT88), .B1(new_n740), .B2(G16), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n741), .B(new_n742), .C1(new_n556), .C2(new_n704), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1341), .ZN(new_n744));
  NOR2_X1   g319(.A1(G171), .A2(new_n704), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G5), .B2(new_n704), .ZN(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n725), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n725), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT29), .B(G2090), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n704), .A2(G4), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n623), .B2(new_n704), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n753), .B(new_n757), .C1(new_n747), .C2(new_n746), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n485), .A2(G103), .A3(G2104), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT25), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n483), .A2(G139), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n485), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n725), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n725), .B2(G33), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT90), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n766), .A2(KEYINPUT90), .A3(new_n767), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n744), .B(new_n758), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n725), .A2(G32), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G141), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT91), .Z(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n479), .A2(G105), .ZN(new_n777));
  INV_X1    g352(.A(G129), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n640), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n771), .B1(new_n780), .B2(new_n725), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT27), .ZN(new_n782));
  INV_X1    g357(.A(G1996), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n725), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n471), .A2(new_n465), .A3(G128), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT89), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n483), .A2(G140), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n485), .A2(G116), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n786), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT31), .B(G11), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT30), .B(G28), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n725), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NOR2_X1   g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n481), .A2(G29), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G2084), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n797), .B1(new_n725), .B2(new_n641), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n766), .B2(new_n767), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n704), .A2(G21), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G168), .B2(new_n704), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n801), .A2(new_n802), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n794), .A2(new_n804), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n784), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n704), .A2(G20), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT23), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n620), .B2(new_n704), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1956), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n725), .A2(G27), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G164), .B2(new_n725), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2078), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n770), .A2(new_n812), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n739), .A2(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NAND2_X1  g399(.A1(new_n623), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n514), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n505), .B1(new_n829), .B2(KEYINPUT95), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT95), .B2(new_n829), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n529), .A2(G55), .B1(G93), .B2(new_n541), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n555), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n555), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n826), .B(new_n836), .Z(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  INV_X1    g418(.A(new_n780), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n497), .A2(new_n499), .ZN(new_n845));
  INV_X1    g420(.A(new_n495), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n792), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n764), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n792), .A2(new_n847), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n849), .B1(new_n848), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n844), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n792), .B(new_n847), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n764), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n780), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n733), .B(new_n632), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n471), .A2(new_n465), .A3(G130), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT96), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n483), .A2(G142), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n485), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n859), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT97), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n854), .A2(new_n866), .A3(new_n857), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT98), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n854), .A2(new_n866), .A3(new_n872), .A4(new_n857), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n866), .B1(new_n854), .B2(new_n857), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n869), .A2(new_n871), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n641), .B(new_n481), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n488), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n882), .B2(new_n868), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT40), .B1(new_n880), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(G395));
  NAND2_X1  g461(.A1(new_n833), .A2(new_n614), .ZN(new_n887));
  NAND2_X1  g462(.A1(G299), .A2(new_n613), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(G299), .A2(new_n613), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT41), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n835), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n555), .A2(new_n833), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n628), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n834), .A2(new_n627), .A3(new_n835), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n892), .A2(new_n888), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(KEYINPUT99), .A3(KEYINPUT41), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n896), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n903), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(new_n900), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G290), .B(G288), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(new_n715), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G290), .B(new_n706), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT101), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n911), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n896), .A2(new_n901), .A3(new_n904), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT100), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n908), .A2(new_n919), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n908), .A2(new_n919), .A3(new_n922), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT102), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n917), .B(KEYINPUT42), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n921), .A2(KEYINPUT100), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n905), .A2(new_n907), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n926), .B(KEYINPUT103), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n923), .A2(new_n925), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n887), .B1(new_n933), .B2(new_n614), .ZN(G295));
  OAI21_X1  g509(.A(new_n887), .B1(new_n933), .B2(new_n614), .ZN(G331));
  XOR2_X1   g510(.A(G286), .B(G301), .Z(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n836), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n834), .A2(new_n835), .A3(new_n936), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n906), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n939), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(KEYINPUT104), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n836), .A2(new_n943), .A3(new_n937), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n896), .A2(new_n904), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n917), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT105), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI221_X1 g525(.A(new_n940), .B1(new_n948), .B2(KEYINPUT105), .C1(new_n945), .C2(new_n946), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT43), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n906), .A2(new_n939), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n942), .B2(new_n944), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n938), .A2(new_n939), .B1(new_n891), .B2(new_n894), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n917), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n956), .B(new_n957), .C1(new_n947), .C2(new_n917), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n952), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n950), .B2(new_n951), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(G397));
  NOR2_X1   g541(.A1(new_n500), .A2(G1384), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n479), .A2(G101), .ZN(new_n969));
  INV_X1    g544(.A(G137), .ZN(new_n970));
  OAI211_X1 g545(.A(G40), .B(new_n969), .C1(new_n477), .C2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n468), .B2(new_n471), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1996), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n780), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n792), .B(G2067), .Z(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n783), .B2(new_n780), .ZN(new_n979));
  INV_X1    g554(.A(new_n973), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n733), .B(new_n736), .Z(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT48), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n734), .A2(new_n736), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT126), .Z(new_n989));
  NOR2_X1   g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n792), .A2(G2067), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n980), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n976), .B(new_n994), .Z(new_n995));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n973), .B1(new_n978), .B2(new_n780), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(KEYINPUT127), .B2(new_n993), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n995), .B2(new_n998), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n987), .B(new_n992), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n972), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n847), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT45), .B(new_n1005), .C1(new_n501), .C2(new_n503), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n807), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1004), .B1(new_n967), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT113), .B(G2084), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n847), .A2(new_n502), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1014), .C1(new_n1017), .C2(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1011), .A2(G168), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(G168), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT51), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1023), .A3(G8), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n578), .A2(new_n586), .A3(G8), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT108), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(KEYINPUT108), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1005), .B1(new_n501), .B2(new_n503), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT50), .ZN(new_n1037));
  INV_X1    g612(.A(G2090), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1013), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT107), .B(G1971), .Z(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1007), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1004), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1035), .B(G8), .C1(new_n1039), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n967), .A2(new_n972), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(new_n709), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n709), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(G8), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1050), .B(new_n1046), .C1(new_n967), .C2(new_n972), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1045), .A2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n1055));
  NOR3_X1   g630(.A1(G305), .A2(new_n1055), .A3(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT109), .B1(new_n715), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT110), .B1(new_n715), .B2(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n1061));
  NAND3_X1  g636(.A1(G305), .A2(new_n1061), .A3(G1981), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT111), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1054), .B1(new_n1064), .B2(KEYINPUT49), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT111), .B(new_n1066), .C1(new_n1059), .C2(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1053), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1042), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1040), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n972), .B1(new_n967), .B2(new_n1012), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1012), .B(new_n1005), .C1(new_n501), .C2(new_n503), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT112), .B(new_n972), .C1(new_n967), .C2(new_n1012), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1074), .A2(new_n1038), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1050), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1044), .B(new_n1068), .C1(new_n1078), .C2(new_n1035), .ZN(new_n1079));
  INV_X1    g654(.A(G2078), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1008), .A2(new_n1009), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT121), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1008), .A2(new_n1009), .A3(new_n1083), .A4(new_n1080), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(KEYINPUT53), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1080), .B(new_n1042), .C1(new_n1017), .C2(KEYINPUT45), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1013), .B1(new_n1017), .B2(new_n1012), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT122), .B(G1961), .Z(new_n1089));
  AOI22_X1  g664(.A1(new_n1086), .A2(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1079), .A2(G301), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1026), .A2(new_n1028), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G288), .A2(G1976), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1059), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1068), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1096), .A2(new_n1054), .B1(new_n1097), .B2(new_n1044), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G168), .A2(G8), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1079), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1100), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1044), .A4(new_n1068), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1098), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1093), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT116), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1042), .B(new_n1112), .C1(new_n1017), .C2(KEYINPUT45), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1041), .A2(new_n1115), .A3(new_n1042), .A4(new_n1112), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT114), .B(G1956), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1114), .A2(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n575), .B2(KEYINPUT115), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G299), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n570), .B(new_n575), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1110), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1123), .B(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1129), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1045), .A2(G2067), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1088), .B2(new_n756), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n623), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1041), .A2(new_n783), .A3(new_n1042), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(G1341), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1045), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1137), .B1(new_n1142), .B2(new_n556), .ZN(new_n1143));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n555), .C1(new_n1138), .C2(new_n1141), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1136), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n972), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(KEYINPUT50), .B2(new_n1036), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1147), .A2(G1348), .B1(G2067), .B2(new_n1045), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n623), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1134), .A2(new_n613), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1135), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1129), .A2(new_n1130), .A3(new_n1123), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1110), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1132), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1149), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1154), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n1160));
  AOI21_X1  g735(.A(G301), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n468), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n485), .B1(new_n468), .B2(new_n1164), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n971), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT124), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1087), .B(G2078), .C1(new_n967), .C2(KEYINPUT45), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1167), .B(new_n1171), .C1(KEYINPUT45), .C2(new_n967), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AND4_X1   g748(.A1(G301), .A2(new_n1162), .A3(new_n1163), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1160), .B1(new_n1161), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1162), .A2(new_n1163), .A3(new_n1173), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(G171), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1085), .A2(new_n1090), .A3(G301), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(KEYINPUT54), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1044), .A2(new_n1068), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1035), .B1(new_n1181), .B2(G8), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1025), .A2(new_n1175), .A3(new_n1179), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1156), .A2(new_n1159), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1109), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(G290), .B(G1986), .Z(new_n1189));
  OAI21_X1  g764(.A(new_n984), .B1(new_n973), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1003), .B1(new_n1188), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g766(.A1(new_n963), .A2(new_n964), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G227), .A2(new_n462), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n702), .A2(new_n661), .A3(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g769(.A(new_n874), .B(KEYINPUT97), .ZN(new_n1196));
  AND2_X1   g770(.A1(new_n871), .A2(new_n873), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n881), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(new_n883), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g774(.A1(new_n1193), .A2(new_n1200), .ZN(G308));
  OAI221_X1 g775(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .C1(new_n963), .C2(new_n964), .ZN(G225));
endmodule


