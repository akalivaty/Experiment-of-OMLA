//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G110), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT24), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n197), .B2(new_n199), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n193), .B2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n205), .A2(new_n206), .A3(new_n194), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n196), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n203), .A2(new_n208), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(KEYINPUT75), .A3(G125), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(KEYINPUT16), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n207), .A2(KEYINPUT74), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n206), .A3(new_n194), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n196), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n201), .A2(new_n202), .ZN(new_n231));
  INV_X1    g045(.A(new_n195), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n198), .A2(G110), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n196), .A2(KEYINPUT24), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT72), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n236), .A2(new_n232), .A3(new_n230), .A4(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n229), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n219), .A2(new_n209), .A3(new_n221), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n209), .B1(new_n219), .B2(new_n221), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n224), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G137), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n245), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n236), .A2(new_n232), .A3(new_n237), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT73), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n251), .A2(new_n238), .B1(new_n228), .B2(new_n225), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n219), .A2(new_n209), .A3(new_n221), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n223), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n248), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n224), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n249), .A2(new_n188), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n257), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n190), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n249), .A2(new_n257), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n189), .A2(G902), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT76), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  OR2_X1    g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT64), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n209), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n271), .A4(new_n270), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT11), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(G137), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(G137), .ZN(new_n285));
  INV_X1    g099(.A(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT11), .A3(G134), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n284), .A2(new_n287), .A3(new_n290), .A4(new_n285), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT65), .B1(new_n278), .B2(new_n271), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n273), .A2(new_n294), .A3(KEYINPUT0), .A4(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n281), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n273), .A2(new_n298), .A3(G128), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n191), .B1(new_n275), .B2(KEYINPUT1), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n273), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n283), .A2(G137), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n286), .A2(G134), .ZN(new_n303));
  OAI21_X1  g117(.A(G131), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n291), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n193), .A2(G116), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT2), .B(G113), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n297), .A2(new_n313), .A3(new_n306), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n269), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n269), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n322), .A2(new_n246), .A3(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n297), .A2(new_n313), .A3(new_n306), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT69), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n316), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT66), .B(KEYINPUT30), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n297), .A2(new_n306), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT30), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n297), .B2(new_n306), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT67), .B(new_n314), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n297), .A2(new_n306), .A3(new_n334), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n280), .A2(new_n274), .B1(new_n293), .B2(new_n295), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n342), .A2(new_n292), .B1(new_n301), .B2(new_n305), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n343), .B2(new_n337), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT67), .B1(new_n344), .B2(new_n314), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n333), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT31), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n333), .B(KEYINPUT31), .C1(new_n340), .C2(new_n345), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n327), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(G472), .A2(G902), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT70), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n327), .ZN(new_n354));
  INV_X1    g168(.A(new_n349), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n314), .B1(new_n335), .B2(new_n338), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n339), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT31), .B1(new_n359), .B2(new_n333), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n354), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n351), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT32), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n348), .A2(new_n349), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n352), .B1(new_n366), .B2(new_n354), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n313), .B1(new_n297), .B2(new_n306), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT28), .B1(new_n329), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT71), .B1(new_n369), .B2(new_n318), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT71), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n317), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n320), .B2(new_n326), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n329), .B1(new_n358), .B2(new_n339), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n326), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n367), .A2(KEYINPUT32), .B1(G472), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n268), .B1(new_n365), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n383));
  NOR2_X1   g197(.A1(G475), .A2(G902), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n322), .A2(new_n246), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n276), .A2(KEYINPUT91), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT91), .B(G143), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT17), .A3(G131), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n385), .A2(new_n386), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n388), .A2(new_n385), .ZN(new_n392));
  OAI21_X1  g206(.A(G131), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n387), .B(new_n290), .C1(new_n385), .C2(new_n388), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n243), .B(new_n390), .C1(KEYINPUT17), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n214), .A2(new_n209), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n217), .A2(new_n218), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(new_n209), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT18), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(new_n290), .ZN(new_n401));
  OAI221_X1 g215(.A(new_n399), .B1(new_n389), .B2(new_n401), .C1(new_n393), .C2(new_n400), .ZN(new_n402));
  XNOR2_X1  g216(.A(G113), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT92), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n396), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n214), .A2(KEYINPUT19), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n398), .B2(KEYINPUT19), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n395), .B(new_n223), .C1(G146), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n410), .B2(new_n402), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n383), .B(new_n384), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT93), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n402), .ZN(new_n414));
  INV_X1    g228(.A(new_n405), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n396), .A2(new_n402), .A3(new_n406), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n384), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT20), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT93), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n418), .A2(new_n421), .A3(new_n383), .A4(new_n384), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n405), .B1(new_n396), .B2(new_n402), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n188), .B1(new_n407), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G475), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT95), .B(G952), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(G234), .A2(G237), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(G898), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(G902), .A3(G953), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n309), .A3(G122), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G122), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT14), .B1(new_n441), .B2(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(G116), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n442), .A2(new_n438), .A3(new_n439), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n444), .A3(G107), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n309), .A2(G122), .ZN(new_n447));
  INV_X1    g261(.A(G107), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n276), .A2(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n191), .A2(G143), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n283), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n283), .B1(new_n451), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n443), .B2(new_n447), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n453), .B1(new_n449), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n276), .A2(G128), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n451), .ZN(new_n461));
  INV_X1    g275(.A(new_n451), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT13), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n283), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  OAI22_X1  g278(.A1(new_n446), .A2(new_n456), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(G217), .A3(new_n246), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OAI221_X1 g284(.A(new_n468), .B1(new_n464), .B2(new_n458), .C1(new_n446), .C2(new_n456), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n188), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(G478), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n472), .B(new_n188), .C1(KEYINPUT15), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n427), .A2(new_n436), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n382), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(G221), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n467), .B2(new_n188), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT77), .Z(new_n484));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT12), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n404), .A2(KEYINPUT78), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G104), .ZN(new_n489));
  AOI21_X1  g303(.A(G107), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n448), .A2(G104), .ZN(new_n491));
  OAI21_X1  g305(.A(G101), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n448), .A3(G104), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n490), .B2(new_n493), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n489), .A3(G107), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n492), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n299), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n300), .A2(new_n273), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT80), .B(KEYINPUT1), .C1(new_n276), .C2(G146), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G128), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT80), .B1(new_n275), .B2(KEYINPUT1), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n278), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n299), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT78), .B(G104), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT3), .B1(new_n509), .B2(G107), .ZN(new_n510));
  AOI21_X1  g324(.A(G101), .B1(new_n509), .B2(G107), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n494), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n512), .A3(new_n492), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n486), .B1(new_n514), .B2(new_n292), .ZN(new_n515));
  INV_X1    g329(.A(new_n292), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n517));
  AOI211_X1 g331(.A(new_n516), .B(new_n517), .C1(new_n503), .C2(new_n513), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n496), .B(new_n494), .C1(new_n490), .C2(new_n493), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n510), .A2(KEYINPUT79), .A3(new_n496), .A4(new_n494), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(G101), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n522), .A2(new_n527), .A3(G101), .A4(new_n523), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n528), .A3(new_n342), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT10), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n513), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n499), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n502), .A2(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n512), .A2(KEYINPUT81), .A3(new_n492), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n529), .A2(new_n516), .A3(new_n531), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G140), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n246), .A2(G227), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n519), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n528), .A2(new_n342), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n497), .B1(new_n520), .B2(new_n521), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n523), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n531), .B(new_n536), .C1(new_n543), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n292), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n541), .B1(new_n548), .B2(new_n537), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n519), .A2(new_n537), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT83), .A3(new_n541), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G469), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n188), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n537), .A3(new_n541), .ZN(new_n557));
  OAI211_X1 g371(.A(G469), .B(new_n557), .C1(new_n552), .C2(new_n541), .ZN(new_n558));
  NAND2_X1  g372(.A1(G469), .A2(G902), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n484), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G110), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT86), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT8), .Z(new_n565));
  INV_X1    g379(.A(G113), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n309), .A2(G119), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT5), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT5), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(KEYINPUT84), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT84), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n311), .A2(new_n312), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n499), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n570), .B2(new_n569), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n565), .B(new_n575), .C1(new_n499), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n502), .A2(new_n212), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n212), .B2(new_n342), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n246), .A2(G224), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT87), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT7), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n582), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n526), .A2(new_n314), .A3(new_n528), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n533), .A2(new_n535), .A3(new_n574), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n564), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n533), .A2(KEYINPUT85), .A3(new_n574), .A4(new_n535), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n586), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n564), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT6), .A3(new_n592), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT6), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n598), .A3(new_n564), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n579), .B(new_n581), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT88), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n597), .A2(KEYINPUT88), .A3(new_n599), .A4(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n594), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G210), .B1(G237), .B2(G902), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT90), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(KEYINPUT89), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n594), .B(new_n609), .C1(new_n603), .C2(new_n604), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n481), .B(new_n562), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n480), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n497), .ZN(G3));
  INV_X1    g429(.A(new_n481), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n603), .A2(new_n604), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n593), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n618), .B2(new_n608), .ZN(new_n619));
  INV_X1    g433(.A(new_n436), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n472), .A2(KEYINPUT96), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n470), .A2(new_n471), .A3(new_n621), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n465), .A2(KEYINPUT97), .A3(new_n468), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n465), .A2(KEYINPUT97), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n621), .B1(new_n627), .B2(new_n469), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n622), .A2(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n476), .A2(G902), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n629), .A2(new_n630), .B1(new_n476), .B2(new_n473), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n423), .B2(new_n426), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n594), .B(new_n608), .C1(new_n603), .C2(new_n604), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n619), .A2(new_n620), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n350), .B2(G902), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n262), .A2(new_n267), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n353), .A2(new_n636), .A3(new_n363), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n484), .ZN(new_n639));
  AOI211_X1 g453(.A(G469), .B(G902), .C1(new_n551), .C2(new_n553), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n639), .B1(new_n640), .B2(new_n560), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  OAI21_X1  g460(.A(new_n481), .B1(new_n605), .B2(new_n607), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n436), .A3(new_n633), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n418), .A2(new_n383), .A3(new_n384), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n383), .B1(new_n418), .B2(new_n384), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n478), .B(new_n426), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n643), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT35), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n248), .A2(KEYINPUT36), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI221_X4 g472(.A(KEYINPUT98), .B1(new_n215), .B2(new_n223), .C1(new_n252), .C2(new_n254), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n255), .B2(new_n224), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n658), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n244), .A2(KEYINPUT98), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n255), .A2(new_n660), .A3(new_n224), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n657), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n266), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n260), .A2(new_n261), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n189), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n479), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n353), .A2(new_n636), .A3(new_n363), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n613), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT37), .B(G110), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR2_X1   g489(.A1(new_n647), .A2(new_n633), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n434), .A2(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n431), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n651), .B2(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n420), .A2(new_n412), .B1(G475), .B2(new_n425), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(KEYINPUT99), .A3(new_n478), .A4(new_n679), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n683), .A3(new_n669), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n365), .B2(new_n381), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n676), .A2(new_n685), .A3(new_n562), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  OAI21_X1  g501(.A(new_n328), .B1(new_n329), .B2(new_n368), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n346), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n188), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n367), .A2(KEYINPUT32), .B1(G472), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n365), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n478), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n423), .B2(new_n426), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(new_n481), .A3(new_n668), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n679), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n562), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n695), .B1(KEYINPUT40), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n611), .A2(new_n612), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT38), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n618), .A2(new_n609), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n605), .A2(new_n610), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT38), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NAND3_X1  g522(.A1(new_n632), .A2(new_n669), .A3(new_n679), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n365), .B2(new_n381), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n619), .A2(new_n562), .A3(new_n634), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT100), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n647), .A2(new_n641), .A3(new_n633), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n710), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  AOI21_X1  g532(.A(new_n555), .B1(new_n554), .B2(new_n188), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n719), .A2(new_n640), .A3(new_n483), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n382), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n635), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NOR2_X1   g538(.A1(new_n653), .A2(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n309), .ZN(G18));
  NAND2_X1  g540(.A1(new_n365), .A2(new_n381), .ZN(new_n727));
  INV_X1    g541(.A(new_n670), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n676), .A2(new_n727), .A3(new_n728), .A4(new_n720), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AND2_X1   g544(.A1(new_n694), .A2(new_n620), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n268), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n637), .A2(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n371), .B1(new_n317), .B2(new_n319), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n369), .A2(KEYINPUT71), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n326), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n348), .B2(new_n349), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT101), .B1(new_n739), .B2(new_n352), .ZN(new_n740));
  INV_X1    g554(.A(new_n738), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n355), .B2(new_n360), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT101), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n351), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n636), .A2(new_n731), .A3(new_n735), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n676), .A3(new_n720), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AOI211_X1 g562(.A(new_n680), .B(new_n631), .C1(new_n426), .C2(new_n423), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n745), .A2(new_n749), .A3(new_n636), .A4(new_n669), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n676), .A3(new_n720), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  AOI21_X1  g567(.A(new_n483), .B1(new_n556), .B2(new_n561), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n702), .A2(new_n481), .A3(new_n703), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n367), .A2(KEYINPUT32), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n380), .A2(G472), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n364), .B1(new_n350), .B2(new_n352), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n749), .A3(new_n735), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT42), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n762));
  INV_X1    g576(.A(new_n749), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(KEYINPUT42), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n382), .A3(new_n764), .A4(new_n754), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n290), .ZN(G33));
  AND2_X1   g581(.A1(new_n681), .A2(new_n683), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n382), .A3(new_n768), .A4(new_n754), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT103), .B(G134), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G36));
  INV_X1    g585(.A(new_n762), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n671), .A2(new_n669), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n629), .A2(new_n630), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n473), .A2(new_n476), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n423), .A3(new_n426), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n777), .A2(new_n423), .A3(KEYINPUT43), .A4(new_n426), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT106), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT107), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n774), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n772), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n557), .B1(new_n552), .B2(new_n541), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT45), .B(new_n557), .C1(new_n552), .C2(new_n541), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n559), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n559), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n556), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n483), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n800), .A3(new_n696), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT104), .ZN(new_n802));
  OAI211_X1 g616(.A(KEYINPUT44), .B(new_n774), .C1(new_n785), .C2(new_n786), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n789), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NOR4_X1   g619(.A1(new_n772), .A2(new_n727), .A3(new_n637), .A4(new_n763), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n800), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n799), .A2(KEYINPUT47), .A3(new_n800), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT108), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT108), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  INV_X1    g632(.A(new_n720), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n772), .A2(new_n431), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n745), .A2(new_n636), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n782), .A2(new_n784), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n820), .A2(new_n669), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n692), .A2(new_n268), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n423), .A2(new_n426), .A3(new_n631), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n821), .A2(new_n735), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n828), .A2(new_n432), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(new_n822), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n706), .A2(new_n701), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n819), .A2(new_n481), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(KEYINPUT115), .A3(new_n832), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n827), .B1(new_n835), .B2(KEYINPUT50), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n830), .B(new_n837), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n432), .A2(new_n828), .A3(new_n822), .A4(new_n762), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n719), .A2(new_n640), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n484), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n809), .A2(new_n844), .A3(new_n810), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n818), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n846), .B2(KEYINPUT51), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n836), .A2(new_n838), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n820), .A2(new_n632), .A3(new_n824), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n829), .A2(new_n822), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n676), .A2(new_n720), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n851), .B(new_n429), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n759), .A2(new_n735), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n820), .A2(new_n855), .A3(new_n822), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n715), .A2(new_n676), .A3(new_n562), .A4(new_n710), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n715), .B1(new_n714), .B2(new_n710), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n679), .B(KEYINPUT112), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT113), .B1(new_n668), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n869));
  INV_X1    g683(.A(new_n867), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n262), .A2(new_n666), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n365), .B2(new_n691), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n676), .A2(new_n873), .A3(new_n694), .A4(new_n754), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n752), .A2(new_n874), .A3(new_n686), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n865), .A2(new_n866), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n752), .A2(new_n874), .A3(new_n686), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(new_n877), .B2(new_n717), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n613), .B1(new_n480), .B2(new_n672), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n725), .A2(new_n880), .A3(new_n722), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n427), .A2(new_n478), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n777), .B1(new_n426), .B2(new_n423), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n436), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n642), .A2(new_n704), .A3(new_n481), .A4(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n747), .A2(new_n729), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n761), .A2(new_n765), .A3(new_n769), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT111), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n751), .A2(new_n762), .A3(new_n888), .A4(new_n754), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT111), .B1(new_n755), .B2(new_n750), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n478), .A2(new_n680), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n682), .A2(KEYINPUT110), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT110), .B1(new_n682), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n668), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n562), .A2(new_n727), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n889), .A2(new_n890), .B1(new_n895), .B2(new_n762), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n881), .A2(new_n886), .A3(new_n887), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n862), .B1(new_n879), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n880), .A2(new_n722), .ZN(new_n899));
  INV_X1    g713(.A(new_n725), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n886), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n887), .A2(new_n896), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n866), .B1(new_n865), .B2(new_n875), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n877), .A2(new_n717), .A3(KEYINPUT52), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n906), .A3(KEYINPUT53), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n898), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n861), .A2(new_n912), .B1(G952), .B2(G953), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n843), .B(KEYINPUT49), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n735), .A2(new_n481), .A3(new_n639), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n915), .A2(new_n692), .A3(new_n778), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n831), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n917), .ZN(G75));
  NOR3_X1   g732(.A1(new_n879), .A2(new_n862), .A3(new_n897), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n903), .B2(new_n906), .ZN(new_n920));
  OAI211_X1 g734(.A(G902), .B(new_n607), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n597), .A2(new_n599), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n600), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n923), .B(new_n924), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n921), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n246), .A2(G952), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT120), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n188), .B1(new_n898), .B2(new_n907), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n932), .B2(new_n607), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT118), .B1(new_n933), .B2(new_n926), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n921), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n937), .A3(new_n925), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n931), .B1(new_n934), .B2(new_n938), .ZN(G51));
  XOR2_X1   g753(.A(new_n559), .B(KEYINPUT57), .Z(new_n940));
  AND3_X1   g754(.A1(new_n898), .A2(new_n907), .A3(new_n910), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n910), .B1(new_n898), .B2(new_n907), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n554), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n794), .B(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n932), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n929), .B1(new_n944), .B2(new_n946), .ZN(G54));
  AND2_X1   g761(.A1(KEYINPUT58), .A2(G475), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n932), .A2(new_n418), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n418), .B1(new_n932), .B2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n929), .ZN(G60));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT59), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n629), .B(new_n953), .C1(new_n941), .C2(new_n942), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n930), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n629), .B1(new_n912), .B2(new_n953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(new_n662), .A2(new_n665), .ZN(new_n958));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n958), .B(new_n961), .C1(new_n919), .C2(new_n920), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n898), .B2(new_n907), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n962), .B(new_n930), .C1(new_n263), .C2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  OAI211_X1 g779(.A(KEYINPUT122), .B(new_n930), .C1(new_n963), .C2(new_n263), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n930), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n919), .B2(new_n920), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n264), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n970), .B(new_n962), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(G66));
  INV_X1    g786(.A(G224), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n433), .A2(new_n973), .A3(new_n246), .ZN(new_n974));
  INV_X1    g788(.A(new_n901), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n246), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n922), .B1(G898), .B2(new_n246), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  AOI21_X1  g792(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n344), .B(new_n409), .Z(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n717), .A2(new_n686), .A3(new_n752), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n707), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n707), .A3(KEYINPUT62), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n562), .A2(new_n696), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n882), .A2(new_n883), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n762), .A2(new_n991), .A3(new_n382), .A4(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n804), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n804), .B2(new_n993), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n989), .B(new_n816), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n983), .B1(new_n996), .B2(new_n246), .ZN(new_n997));
  INV_X1    g811(.A(new_n982), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n802), .A2(new_n676), .A3(new_n694), .A4(new_n855), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n887), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n804), .A3(new_n816), .A4(new_n984), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n979), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n979), .ZN(new_n1006));
  INV_X1    g820(.A(new_n995), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n804), .A2(new_n990), .A3(new_n993), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g823(.A1(new_n987), .A2(new_n988), .B1(new_n815), .B2(new_n813), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1006), .B(new_n1003), .C1(new_n1011), .C2(new_n983), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1005), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n1002), .B2(new_n901), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n378), .A2(new_n328), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n346), .B1(new_n378), .B2(new_n326), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n908), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1019), .B(new_n1021), .C1(G952), .C2(new_n246), .ZN(new_n1022));
  INV_X1    g836(.A(new_n378), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n326), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1009), .A2(new_n1010), .A3(new_n975), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(new_n1015), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1022), .A2(new_n1026), .ZN(G57));
endmodule


