

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743;

  INV_X1 U368 ( .A(G953), .ZN(n719) );
  XNOR2_X2 U369 ( .A(n575), .B(n574), .ZN(n600) );
  INV_X2 U370 ( .A(n654), .ZN(n594) );
  NOR2_X1 U371 ( .A1(n667), .A2(n591), .ZN(n352) );
  XNOR2_X1 U372 ( .A(G131), .B(G134), .ZN(n441) );
  XNOR2_X1 U373 ( .A(n352), .B(KEYINPUT34), .ZN(n567) );
  XNOR2_X1 U374 ( .A(n450), .B(n449), .ZN(n545) );
  OR2_X2 U375 ( .A1(n710), .A2(G902), .ZN(n382) );
  XNOR2_X1 U376 ( .A(n468), .B(n348), .ZN(n381) );
  XNOR2_X1 U377 ( .A(n441), .B(KEYINPUT66), .ZN(n483) );
  XNOR2_X2 U378 ( .A(n577), .B(n365), .ZN(n392) );
  XNOR2_X2 U379 ( .A(n582), .B(n349), .ZN(n393) );
  XNOR2_X1 U380 ( .A(n538), .B(KEYINPUT86), .ZN(n373) );
  NAND2_X1 U381 ( .A1(n696), .A2(n539), .ZN(n372) );
  XNOR2_X1 U382 ( .A(n501), .B(n429), .ZN(n455) );
  XNOR2_X1 U383 ( .A(G140), .B(KEYINPUT10), .ZN(n429) );
  XNOR2_X1 U384 ( .A(n545), .B(KEYINPUT1), .ZN(n556) );
  INV_X1 U385 ( .A(G472), .ZN(n412) );
  INV_X1 U386 ( .A(KEYINPUT91), .ZN(n404) );
  OR2_X1 U387 ( .A1(n742), .A2(n603), .ZN(n583) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n481) );
  INV_X2 U389 ( .A(G146), .ZN(n446) );
  INV_X1 U390 ( .A(G237), .ZN(n488) );
  XNOR2_X1 U391 ( .A(n453), .B(KEYINPUT21), .ZN(n643) );
  NOR2_X1 U392 ( .A1(n380), .A2(n697), .ZN(n379) );
  NOR2_X1 U393 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U394 ( .A(n445), .B(KEYINPUT4), .ZN(n729) );
  XNOR2_X1 U395 ( .A(n394), .B(G107), .ZN(n495) );
  INV_X1 U396 ( .A(G116), .ZN(n394) );
  XOR2_X1 U397 ( .A(G104), .B(G107), .Z(n443) );
  XNOR2_X1 U398 ( .A(n729), .B(G101), .ZN(n497) );
  XNOR2_X1 U399 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n499) );
  NOR2_X1 U400 ( .A1(n628), .A2(n346), .ZN(n411) );
  XNOR2_X1 U401 ( .A(n361), .B(n360), .ZN(n714) );
  XNOR2_X1 U402 ( .A(n362), .B(n496), .ZN(n361) );
  XNOR2_X1 U403 ( .A(n494), .B(n493), .ZN(n360) );
  XNOR2_X1 U404 ( .A(n495), .B(KEYINPUT16), .ZN(n362) );
  XNOR2_X1 U405 ( .A(KEYINPUT23), .B(KEYINPUT73), .ZN(n456) );
  XNOR2_X1 U406 ( .A(KEYINPUT94), .B(KEYINPUT15), .ZN(n451) );
  XNOR2_X1 U407 ( .A(n353), .B(n370), .ZN(n667) );
  INV_X1 U408 ( .A(KEYINPUT33), .ZN(n370) );
  XNOR2_X1 U409 ( .A(n506), .B(KEYINPUT90), .ZN(n507) );
  XNOR2_X1 U410 ( .A(n356), .B(KEYINPUT19), .ZN(n563) );
  NOR2_X1 U411 ( .A1(n535), .A2(n357), .ZN(n356) );
  NOR2_X1 U412 ( .A1(n700), .A2(G902), .ZN(n450) );
  XNOR2_X1 U413 ( .A(KEYINPUT108), .B(KEYINPUT28), .ZN(n516) );
  XNOR2_X1 U414 ( .A(n654), .B(KEYINPUT6), .ZN(n598) );
  OR2_X1 U415 ( .A1(n743), .A2(n741), .ZN(n375) );
  OR2_X1 U416 ( .A1(n588), .A2(n403), .ZN(n401) );
  AND2_X1 U417 ( .A1(n584), .A2(n395), .ZN(n402) );
  XOR2_X1 U418 ( .A(G116), .B(G113), .Z(n484) );
  XNOR2_X1 U419 ( .A(n482), .B(n387), .ZN(n386) );
  XNOR2_X1 U420 ( .A(G119), .B(KEYINPUT5), .ZN(n387) );
  XNOR2_X1 U421 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n477) );
  XNOR2_X1 U422 ( .A(G143), .B(G131), .ZN(n433) );
  XNOR2_X1 U423 ( .A(G113), .B(G104), .ZN(n430) );
  BUF_X1 U424 ( .A(n455), .Z(n727) );
  XNOR2_X1 U425 ( .A(n510), .B(KEYINPUT109), .ZN(n637) );
  NOR2_X1 U426 ( .A1(n515), .A2(n514), .ZN(n540) );
  INV_X1 U427 ( .A(G902), .ZN(n489) );
  NOR2_X1 U428 ( .A1(n378), .A2(n376), .ZN(n732) );
  XNOR2_X1 U429 ( .A(G134), .B(G122), .ZN(n419) );
  XOR2_X1 U430 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n421) );
  XNOR2_X1 U431 ( .A(n444), .B(n355), .ZN(n369) );
  XNOR2_X1 U432 ( .A(G140), .B(G110), .ZN(n355) );
  XNOR2_X1 U433 ( .A(n363), .B(n714), .ZN(n622) );
  XNOR2_X1 U434 ( .A(n364), .B(n502), .ZN(n363) );
  NAND2_X1 U435 ( .A1(G237), .A2(G234), .ZN(n471) );
  XNOR2_X1 U436 ( .A(n569), .B(n568), .ZN(n742) );
  XNOR2_X1 U437 ( .A(KEYINPUT35), .B(KEYINPUT82), .ZN(n568) );
  NOR2_X1 U438 ( .A1(n492), .A2(n491), .ZN(n531) );
  AND2_X1 U439 ( .A1(n410), .A2(n408), .ZN(n407) );
  AND2_X1 U440 ( .A1(n409), .A2(n629), .ZN(n408) );
  XNOR2_X1 U441 ( .A(n465), .B(n464), .ZN(n710) );
  AND2_X2 U442 ( .A1(n366), .A2(n358), .ZN(n709) );
  NOR2_X1 U443 ( .A1(n613), .A2(n359), .ZN(n358) );
  INV_X1 U444 ( .A(n612), .ZN(n359) );
  AND2_X1 U445 ( .A1(n671), .A2(n670), .ZN(n672) );
  BUF_X1 U446 ( .A(n742), .Z(n354) );
  NOR2_X1 U447 ( .A1(n656), .A2(n591), .ZN(n592) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n529) );
  INV_X1 U449 ( .A(KEYINPUT84), .ZN(n390) );
  INV_X1 U450 ( .A(KEYINPUT107), .ZN(n365) );
  XNOR2_X1 U451 ( .A(n392), .B(G110), .ZN(G12) );
  INV_X1 U452 ( .A(n671), .ZN(n413) );
  NAND2_X1 U453 ( .A1(n366), .A2(n612), .ZN(n671) );
  OR2_X1 U454 ( .A1(n613), .A2(n412), .ZN(n346) );
  INV_X1 U455 ( .A(n713), .ZN(n629) );
  XNOR2_X1 U456 ( .A(n430), .B(G122), .ZN(n494) );
  OR2_X1 U457 ( .A1(n698), .A2(KEYINPUT88), .ZN(n347) );
  BUF_X1 U458 ( .A(n556), .Z(n648) );
  XOR2_X1 U459 ( .A(n466), .B(KEYINPUT81), .Z(n348) );
  XOR2_X1 U460 ( .A(KEYINPUT83), .B(KEYINPUT32), .Z(n349) );
  XOR2_X1 U461 ( .A(n614), .B(KEYINPUT59), .Z(n350) );
  XOR2_X1 U462 ( .A(n622), .B(n621), .Z(n351) );
  XNOR2_X1 U463 ( .A(n617), .B(KEYINPUT93), .ZN(n713) );
  XNOR2_X1 U464 ( .A(n609), .B(n608), .ZN(n718) );
  NAND2_X1 U465 ( .A1(n602), .A2(n404), .ZN(n403) );
  NAND2_X1 U466 ( .A1(n414), .A2(n598), .ZN(n353) );
  NAND2_X1 U467 ( .A1(n553), .A2(KEYINPUT88), .ZN(n377) );
  NAND2_X1 U468 ( .A1(n718), .A2(n732), .ZN(n367) );
  INV_X1 U469 ( .A(n632), .ZN(n357) );
  XNOR2_X2 U470 ( .A(n505), .B(n504), .ZN(n535) );
  INV_X1 U471 ( .A(n497), .ZN(n364) );
  XNOR2_X2 U472 ( .A(n367), .B(n610), .ZN(n366) );
  XNOR2_X1 U473 ( .A(n476), .B(n368), .ZN(n700) );
  XNOR2_X1 U474 ( .A(n369), .B(n728), .ZN(n368) );
  NAND2_X1 U475 ( .A1(n374), .A2(n371), .ZN(n548) );
  XNOR2_X1 U476 ( .A(n375), .B(n522), .ZN(n374) );
  NAND2_X1 U477 ( .A1(n377), .A2(n379), .ZN(n376) );
  NOR2_X1 U478 ( .A1(n553), .A2(n347), .ZN(n378) );
  AND2_X1 U479 ( .A1(n698), .A2(KEYINPUT88), .ZN(n380) );
  XNOR2_X2 U480 ( .A(n382), .B(n381), .ZN(n579) );
  XNOR2_X1 U481 ( .A(n383), .B(n476), .ZN(n627) );
  XNOR2_X1 U482 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U483 ( .A(n496), .B(n480), .ZN(n384) );
  XNOR2_X1 U484 ( .A(n388), .B(n386), .ZN(n385) );
  XNOR2_X1 U485 ( .A(n483), .B(n484), .ZN(n388) );
  XNOR2_X1 U486 ( .A(n497), .B(n446), .ZN(n476) );
  NAND2_X1 U487 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U488 ( .A1(n519), .A2(n389), .ZN(n391) );
  NOR2_X1 U489 ( .A1(n563), .A2(n545), .ZN(n389) );
  NAND2_X1 U490 ( .A1(n529), .A2(n636), .ZN(n530) );
  NAND2_X1 U491 ( .A1(n392), .A2(n393), .ZN(n603) );
  XNOR2_X1 U492 ( .A(n393), .B(G119), .ZN(G21) );
  NAND2_X1 U493 ( .A1(n584), .A2(KEYINPUT64), .ZN(n405) );
  NOR2_X1 U494 ( .A1(n403), .A2(n585), .ZN(n395) );
  NAND2_X1 U495 ( .A1(n398), .A2(n396), .ZN(n607) );
  NAND2_X1 U496 ( .A1(n405), .A2(n397), .ZN(n396) );
  AND2_X1 U497 ( .A1(n588), .A2(KEYINPUT91), .ZN(n397) );
  NOR2_X1 U498 ( .A1(n402), .A2(n399), .ZN(n398) );
  NAND2_X1 U499 ( .A1(n401), .A2(n400), .ZN(n399) );
  OR2_X1 U500 ( .A1(n602), .A2(n404), .ZN(n400) );
  NAND2_X1 U501 ( .A1(n407), .A2(n406), .ZN(n630) );
  NAND2_X1 U502 ( .A1(n671), .A2(n628), .ZN(n406) );
  NAND2_X1 U503 ( .A1(n628), .A2(n346), .ZN(n409) );
  NAND2_X1 U504 ( .A1(n413), .A2(n411), .ZN(n410) );
  XNOR2_X2 U505 ( .A(G143), .B(G128), .ZN(n445) );
  AND2_X1 U506 ( .A1(n589), .A2(n557), .ZN(n414) );
  XNOR2_X1 U507 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n415) );
  XNOR2_X1 U508 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n416) );
  AND2_X1 U509 ( .A1(n648), .A2(n576), .ZN(n417) );
  AND2_X1 U510 ( .A1(n581), .A2(n580), .ZN(n418) );
  XNOR2_X1 U511 ( .A(n477), .B(KEYINPUT72), .ZN(n496) );
  XNOR2_X1 U512 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT24), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n668), .A2(n527), .ZN(n521) );
  XNOR2_X1 U515 ( .A(n675), .B(n674), .ZN(G75) );
  XNOR2_X1 U516 ( .A(KEYINPUT46), .B(KEYINPUT89), .ZN(n522) );
  XOR2_X1 U517 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n420) );
  XNOR2_X1 U518 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U519 ( .A(n445), .B(n421), .Z(n422) );
  XNOR2_X1 U520 ( .A(n495), .B(n422), .ZN(n423) );
  XOR2_X1 U521 ( .A(n424), .B(n423), .Z(n427) );
  NAND2_X1 U522 ( .A1(G234), .A2(n719), .ZN(n425) );
  XOR2_X1 U523 ( .A(KEYINPUT8), .B(n425), .Z(n461) );
  NAND2_X1 U524 ( .A1(G217), .A2(n461), .ZN(n426) );
  XNOR2_X1 U525 ( .A(n427), .B(n426), .ZN(n706) );
  NOR2_X1 U526 ( .A1(G902), .A2(n706), .ZN(n428) );
  XNOR2_X1 U527 ( .A(G478), .B(n428), .ZN(n523) );
  XNOR2_X2 U528 ( .A(n446), .B(G125), .ZN(n501) );
  XOR2_X1 U529 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n432) );
  NAND2_X1 U530 ( .A1(G214), .A2(n481), .ZN(n431) );
  XNOR2_X1 U531 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n434) );
  XNOR2_X1 U533 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U534 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U535 ( .A(n494), .B(n437), .ZN(n438) );
  XNOR2_X1 U536 ( .A(n727), .B(n438), .ZN(n614) );
  NAND2_X1 U537 ( .A1(n614), .A2(n489), .ZN(n440) );
  XNOR2_X1 U538 ( .A(KEYINPUT13), .B(G475), .ZN(n439) );
  XNOR2_X1 U539 ( .A(n440), .B(n439), .ZN(n524) );
  INV_X1 U540 ( .A(n524), .ZN(n532) );
  NAND2_X1 U541 ( .A1(n523), .A2(n532), .ZN(n690) );
  XNOR2_X1 U542 ( .A(G137), .B(KEYINPUT65), .ZN(n457) );
  XNOR2_X1 U543 ( .A(n483), .B(n457), .ZN(n728) );
  NAND2_X1 U544 ( .A1(G227), .A2(n719), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U546 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n448) );
  INV_X1 U547 ( .A(G469), .ZN(n447) );
  INV_X1 U548 ( .A(n545), .ZN(n518) );
  XNOR2_X1 U549 ( .A(n451), .B(G902), .ZN(n613) );
  NAND2_X1 U550 ( .A1(n613), .A2(G234), .ZN(n452) );
  XNOR2_X1 U551 ( .A(KEYINPUT20), .B(n452), .ZN(n467) );
  NAND2_X1 U552 ( .A1(G221), .A2(n467), .ZN(n453) );
  INV_X1 U553 ( .A(KEYINPUT97), .ZN(n454) );
  XNOR2_X1 U554 ( .A(n643), .B(n454), .ZN(n570) );
  XNOR2_X1 U555 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U556 ( .A(G128), .B(n457), .ZN(n458) );
  XNOR2_X1 U557 ( .A(n460), .B(n459), .ZN(n465) );
  XOR2_X1 U558 ( .A(G119), .B(G110), .Z(n493) );
  XOR2_X1 U559 ( .A(n493), .B(KEYINPUT95), .Z(n463) );
  NAND2_X1 U560 ( .A1(G221), .A2(n461), .ZN(n462) );
  XNOR2_X1 U561 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U562 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n466) );
  NAND2_X1 U563 ( .A1(G217), .A2(n467), .ZN(n468) );
  NOR2_X2 U564 ( .A1(n570), .A2(n579), .ZN(n589) );
  NAND2_X1 U565 ( .A1(n518), .A2(n589), .ZN(n593) );
  NOR2_X1 U566 ( .A1(G900), .A2(n719), .ZN(n469) );
  NAND2_X1 U567 ( .A1(n469), .A2(G902), .ZN(n470) );
  NAND2_X1 U568 ( .A1(n719), .A2(G952), .ZN(n558) );
  NAND2_X1 U569 ( .A1(n470), .A2(n558), .ZN(n473) );
  XNOR2_X1 U570 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n472), .B(n471), .ZN(n665) );
  INV_X1 U572 ( .A(n665), .ZN(n560) );
  NAND2_X1 U573 ( .A1(n473), .A2(n560), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n593), .A2(n512), .ZN(n475) );
  INV_X1 U575 ( .A(KEYINPUT80), .ZN(n474) );
  XNOR2_X1 U576 ( .A(n475), .B(n474), .ZN(n492) );
  XOR2_X1 U577 ( .A(G137), .B(KEYINPUT78), .Z(n479) );
  XNOR2_X1 U578 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n478) );
  XNOR2_X1 U579 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U580 ( .A1(n481), .A2(G210), .ZN(n482) );
  NAND2_X1 U581 ( .A1(n627), .A2(n489), .ZN(n487) );
  INV_X1 U582 ( .A(KEYINPUT100), .ZN(n485) );
  XNOR2_X1 U583 ( .A(n485), .B(G472), .ZN(n486) );
  XNOR2_X2 U584 ( .A(n487), .B(n486), .ZN(n654) );
  NAND2_X1 U585 ( .A1(n489), .A2(n488), .ZN(n503) );
  NAND2_X1 U586 ( .A1(n503), .A2(G214), .ZN(n632) );
  NAND2_X1 U587 ( .A1(n594), .A2(n632), .ZN(n490) );
  XNOR2_X1 U588 ( .A(KEYINPUT30), .B(n490), .ZN(n491) );
  NAND2_X1 U589 ( .A1(n719), .A2(G224), .ZN(n498) );
  XNOR2_X1 U590 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U591 ( .A(n501), .B(n500), .ZN(n502) );
  NAND2_X1 U592 ( .A1(n622), .A2(n613), .ZN(n505) );
  NAND2_X1 U593 ( .A1(n503), .A2(G210), .ZN(n504) );
  XNOR2_X1 U594 ( .A(n535), .B(KEYINPUT38), .ZN(n631) );
  NAND2_X1 U595 ( .A1(n531), .A2(n631), .ZN(n508) );
  XOR2_X1 U596 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n506) );
  XNOR2_X1 U597 ( .A(n508), .B(n507), .ZN(n555) );
  NOR2_X1 U598 ( .A1(n690), .A2(n555), .ZN(n509) );
  XNOR2_X1 U599 ( .A(n509), .B(KEYINPUT40), .ZN(n743) );
  NAND2_X1 U600 ( .A1(n631), .A2(n632), .ZN(n510) );
  AND2_X1 U601 ( .A1(n524), .A2(n523), .ZN(n635) );
  NAND2_X1 U602 ( .A1(n637), .A2(n635), .ZN(n511) );
  XOR2_X1 U603 ( .A(KEYINPUT41), .B(n511), .Z(n668) );
  INV_X1 U604 ( .A(n579), .ZN(n515) );
  NOR2_X1 U605 ( .A1(n643), .A2(n512), .ZN(n513) );
  XOR2_X1 U606 ( .A(KEYINPUT68), .B(n513), .Z(n514) );
  AND2_X1 U607 ( .A1(n594), .A2(n540), .ZN(n517) );
  XNOR2_X1 U608 ( .A(n517), .B(n516), .ZN(n519) );
  XNOR2_X1 U609 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n520) );
  XNOR2_X1 U610 ( .A(n521), .B(n520), .ZN(n741) );
  INV_X1 U611 ( .A(n523), .ZN(n533) );
  NAND2_X1 U612 ( .A1(n524), .A2(n533), .ZN(n693) );
  XOR2_X1 U613 ( .A(KEYINPUT105), .B(n693), .Z(n554) );
  NAND2_X1 U614 ( .A1(n554), .A2(n690), .ZN(n636) );
  INV_X1 U615 ( .A(n636), .ZN(n525) );
  NOR2_X1 U616 ( .A1(KEYINPUT47), .A2(n525), .ZN(n526) );
  XNOR2_X1 U617 ( .A(n526), .B(KEYINPUT76), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n528), .A2(n529), .ZN(n539) );
  NAND2_X1 U619 ( .A1(n530), .A2(KEYINPUT47), .ZN(n537) );
  INV_X1 U620 ( .A(n531), .ZN(n534) );
  NAND2_X1 U621 ( .A1(n533), .A2(n532), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n534), .A2(n565), .ZN(n536) );
  INV_X1 U623 ( .A(n535), .ZN(n551) );
  NAND2_X1 U624 ( .A1(n536), .A2(n551), .ZN(n676) );
  NAND2_X1 U625 ( .A1(n537), .A2(n676), .ZN(n538) );
  INV_X1 U626 ( .A(n690), .ZN(n688) );
  NAND2_X1 U627 ( .A1(n688), .A2(n632), .ZN(n542) );
  NAND2_X1 U628 ( .A1(n540), .A2(n598), .ZN(n541) );
  NOR2_X1 U629 ( .A1(n542), .A2(n541), .ZN(n549) );
  NAND2_X1 U630 ( .A1(n549), .A2(n551), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n543), .B(KEYINPUT36), .ZN(n544) );
  XNOR2_X1 U632 ( .A(KEYINPUT111), .B(n544), .ZN(n546) );
  NAND2_X1 U633 ( .A1(n546), .A2(n557), .ZN(n696) );
  XOR2_X1 U634 ( .A(KEYINPUT67), .B(KEYINPUT48), .Z(n547) );
  XNOR2_X1 U635 ( .A(n548), .B(n547), .ZN(n553) );
  AND2_X1 U636 ( .A1(n648), .A2(n549), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n550), .B(KEYINPUT43), .ZN(n552) );
  NOR2_X1 U638 ( .A1(n552), .A2(n551), .ZN(n698) );
  NOR2_X1 U639 ( .A1(n555), .A2(n554), .ZN(n697) );
  INV_X1 U640 ( .A(n556), .ZN(n557) );
  NOR2_X1 U641 ( .A1(G898), .A2(n719), .ZN(n717) );
  NAND2_X1 U642 ( .A1(n717), .A2(G902), .ZN(n559) );
  NAND2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X2 U645 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X2 U646 ( .A(n564), .B(KEYINPUT0), .ZN(n573) );
  INV_X1 U647 ( .A(n573), .ZN(n591) );
  INV_X1 U648 ( .A(n565), .ZN(n566) );
  NAND2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n569) );
  INV_X1 U650 ( .A(n570), .ZN(n571) );
  AND2_X1 U651 ( .A1(n635), .A2(n571), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U653 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n574) );
  AND2_X1 U654 ( .A1(n654), .A2(n579), .ZN(n576) );
  NAND2_X1 U655 ( .A1(n600), .A2(n417), .ZN(n577) );
  INV_X1 U656 ( .A(n598), .ZN(n581) );
  INV_X1 U657 ( .A(KEYINPUT106), .ZN(n578) );
  XNOR2_X1 U658 ( .A(n579), .B(n578), .ZN(n642) );
  NOR2_X1 U659 ( .A1(n648), .A2(n642), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n600), .A2(n418), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(KEYINPUT44), .ZN(n584) );
  INV_X1 U662 ( .A(KEYINPUT64), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n585), .A2(KEYINPUT44), .ZN(n586) );
  NOR2_X1 U664 ( .A1(n742), .A2(n586), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n587), .A2(n603), .ZN(n588) );
  INV_X1 U666 ( .A(n589), .ZN(n647) );
  NOR2_X1 U667 ( .A1(n647), .A2(n648), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n590), .A2(n594), .ZN(n656) );
  XNOR2_X1 U669 ( .A(n592), .B(KEYINPUT31), .ZN(n692) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n573), .A2(n595), .ZN(n679) );
  NAND2_X1 U672 ( .A1(n692), .A2(n679), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n596), .A2(n636), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n648), .A2(n642), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n677) );
  AND2_X1 U677 ( .A1(n601), .A2(n677), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n354), .A2(KEYINPUT44), .ZN(n605) );
  XOR2_X1 U679 ( .A(KEYINPUT92), .B(n603), .Z(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT87), .B(KEYINPUT45), .Z(n608) );
  INV_X1 U683 ( .A(KEYINPUT2), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n611), .A2(KEYINPUT79), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(KEYINPUT79), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n709), .A2(G475), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n615), .B(n350), .ZN(n618) );
  INV_X1 U688 ( .A(G952), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n616), .A2(G953), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n629), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n619), .B(n416), .ZN(G60) );
  NAND2_X1 U692 ( .A1(n709), .A2(G210), .ZN(n623) );
  XOR2_X1 U693 ( .A(KEYINPUT85), .B(KEYINPUT54), .Z(n620) );
  XNOR2_X1 U694 ( .A(n620), .B(KEYINPUT55), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n623), .B(n351), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n624), .A2(n629), .ZN(n626) );
  INV_X1 U697 ( .A(KEYINPUT56), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(G51) );
  XOR2_X1 U699 ( .A(KEYINPUT62), .B(n627), .Z(n628) );
  XNOR2_X1 U700 ( .A(n630), .B(n415), .ZN(G57) );
  INV_X1 U701 ( .A(n631), .ZN(n633) );
  NAND2_X1 U702 ( .A1(n633), .A2(n357), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U706 ( .A(KEYINPUT120), .B(n640), .Z(n641) );
  NOR2_X1 U707 ( .A1(n667), .A2(n641), .ZN(n662) );
  INV_X1 U708 ( .A(n642), .ZN(n644) );
  NAND2_X1 U709 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U710 ( .A(n645), .B(KEYINPUT49), .ZN(n646) );
  XNOR2_X1 U711 ( .A(KEYINPUT116), .B(n646), .ZN(n652) );
  NAND2_X1 U712 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U713 ( .A(n649), .B(KEYINPUT117), .ZN(n650) );
  XNOR2_X1 U714 ( .A(KEYINPUT50), .B(n650), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U717 ( .A(n655), .B(KEYINPUT118), .ZN(n657) );
  NAND2_X1 U718 ( .A1(n657), .A2(n656), .ZN(n659) );
  XOR2_X1 U719 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n658) );
  XNOR2_X1 U720 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X1 U721 ( .A1(n660), .A2(n668), .ZN(n661) );
  NOR2_X1 U722 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U723 ( .A(n663), .B(KEYINPUT52), .ZN(n664) );
  NOR2_X1 U724 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U725 ( .A1(n666), .A2(G952), .ZN(n673) );
  NOR2_X1 U726 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U727 ( .A1(n669), .A2(G953), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U729 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n674) );
  XNOR2_X1 U730 ( .A(n676), .B(G143), .ZN(G45) );
  XNOR2_X1 U731 ( .A(G101), .B(n677), .ZN(G3) );
  NOR2_X1 U732 ( .A1(n690), .A2(n679), .ZN(n678) );
  XOR2_X1 U733 ( .A(G104), .B(n678), .Z(G6) );
  NOR2_X1 U734 ( .A1(n679), .A2(n693), .ZN(n683) );
  XOR2_X1 U735 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n681) );
  XNOR2_X1 U736 ( .A(G107), .B(KEYINPUT27), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U738 ( .A(n683), .B(n682), .ZN(G9) );
  XOR2_X1 U739 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n686) );
  INV_X1 U740 ( .A(n693), .ZN(n684) );
  NAND2_X1 U741 ( .A1(n684), .A2(n529), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U743 ( .A(G128), .B(n687), .ZN(G30) );
  NAND2_X1 U744 ( .A1(n529), .A2(n688), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n689), .B(G146), .ZN(G48) );
  NOR2_X1 U746 ( .A1(n690), .A2(n692), .ZN(n691) );
  XOR2_X1 U747 ( .A(G113), .B(n691), .Z(G15) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U749 ( .A(G116), .B(n694), .Z(G18) );
  XOR2_X1 U750 ( .A(G125), .B(KEYINPUT37), .Z(n695) );
  XNOR2_X1 U751 ( .A(n696), .B(n695), .ZN(G27) );
  XOR2_X1 U752 ( .A(G134), .B(n697), .Z(G36) );
  XNOR2_X1 U753 ( .A(n698), .B(G140), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n699), .B(KEYINPUT115), .ZN(G42) );
  XNOR2_X1 U755 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n700), .B(KEYINPUT57), .ZN(n701) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U758 ( .A1(n709), .A2(G469), .ZN(n703) );
  XOR2_X1 U759 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U760 ( .A1(n713), .A2(n705), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n709), .A2(G478), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n713), .A2(n708), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n709), .A2(G217), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(G66) );
  XNOR2_X1 U767 ( .A(n714), .B(G101), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT125), .ZN(n716) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n726) );
  NAND2_X1 U770 ( .A1(n718), .A2(n719), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n720), .B(KEYINPUT124), .ZN(n724) );
  NAND2_X1 U772 ( .A1(G953), .A2(G224), .ZN(n721) );
  XNOR2_X1 U773 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n722), .A2(G898), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(G69) );
  XNOR2_X1 U777 ( .A(n727), .B(KEYINPUT126), .ZN(n731) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U779 ( .A(n731), .B(n730), .Z(n736) );
  BUF_X1 U780 ( .A(n732), .Z(n733) );
  XNOR2_X1 U781 ( .A(n736), .B(n733), .ZN(n734) );
  NOR2_X1 U782 ( .A1(G953), .A2(n734), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n735), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U784 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G953), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(G72) );
  XOR2_X1 U788 ( .A(G137), .B(n741), .Z(G39) );
  XOR2_X1 U789 ( .A(n354), .B(G122), .Z(G24) );
  XOR2_X1 U790 ( .A(n743), .B(G131), .Z(G33) );
endmodule

