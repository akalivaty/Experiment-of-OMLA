

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589;

  AND2_X1 U329 ( .A1(n555), .A2(n532), .ZN(n471) );
  XOR2_X1 U330 ( .A(KEYINPUT28), .B(n469), .Z(n532) );
  XOR2_X1 U331 ( .A(KEYINPUT45), .B(n405), .Z(n297) );
  INV_X1 U332 ( .A(KEYINPUT11), .ZN(n388) );
  XNOR2_X1 U333 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U334 ( .A(n340), .B(n419), .ZN(n341) );
  XNOR2_X1 U335 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U336 ( .A1(n409), .A2(n408), .ZN(n411) );
  XNOR2_X1 U337 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U338 ( .A(n478), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U339 ( .A(n480), .B(n479), .ZN(n525) );
  NOR2_X1 U340 ( .A1(n536), .A2(n451), .ZN(n571) );
  INV_X1 U341 ( .A(G36GAT), .ZN(n484) );
  XNOR2_X1 U342 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U343 ( .A(n484), .B(KEYINPUT106), .ZN(n485) );
  XNOR2_X1 U344 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n486), .B(n485), .ZN(G1329GAT) );
  XOR2_X1 U346 ( .A(G85GAT), .B(G92GAT), .Z(n384) );
  XOR2_X1 U347 ( .A(G57GAT), .B(KEYINPUT13), .Z(n357) );
  XNOR2_X1 U348 ( .A(n384), .B(n357), .ZN(n311) );
  XNOR2_X1 U349 ( .A(G148GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n298), .B(G78GAT), .ZN(n332) );
  XOR2_X1 U351 ( .A(n332), .B(KEYINPUT73), .Z(n300) );
  NAND2_X1 U352 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U354 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n302) );
  XNOR2_X1 U355 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(n304), .B(n303), .Z(n309) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G120GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n305), .B(G71GAT), .ZN(n315) );
  XOR2_X1 U360 ( .A(G204GAT), .B(KEYINPUT72), .Z(n307) );
  XNOR2_X1 U361 ( .A(G176GAT), .B(G64GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n420) );
  XNOR2_X1 U363 ( .A(n315), .B(n420), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n481) );
  XNOR2_X1 U366 ( .A(KEYINPUT41), .B(n481), .ZN(n558) );
  XNOR2_X1 U367 ( .A(KEYINPUT109), .B(n558), .ZN(n540) );
  XOR2_X1 U368 ( .A(KEYINPUT17), .B(G183GAT), .Z(n313) );
  XNOR2_X1 U369 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U371 ( .A(KEYINPUT84), .B(n314), .Z(n424) );
  XOR2_X1 U372 ( .A(n315), .B(G176GAT), .Z(n317) );
  XOR2_X1 U373 ( .A(G190GAT), .B(G134GAT), .Z(n397) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(n397), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n424), .B(n318), .ZN(n327) );
  XOR2_X1 U377 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n320) );
  NAND2_X1 U378 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U380 ( .A(n321), .B(KEYINPUT83), .Z(n325) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G113GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n322), .B(G15GAT), .ZN(n373) );
  XNOR2_X1 U383 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n323), .B(KEYINPUT81), .ZN(n441) );
  XNOR2_X1 U385 ( .A(n373), .B(n441), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n536) );
  XOR2_X1 U388 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n329) );
  XNOR2_X1 U389 ( .A(G50GAT), .B(G204GAT), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n344) );
  XOR2_X1 U391 ( .A(G155GAT), .B(KEYINPUT2), .Z(n331) );
  XNOR2_X1 U392 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n433) );
  XNOR2_X1 U394 ( .A(n433), .B(n332), .ZN(n337) );
  XOR2_X1 U395 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n334) );
  NAND2_X1 U396 ( .A1(G228GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n335), .B(KEYINPUT24), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U400 ( .A(G141GAT), .B(G22GAT), .Z(n377) );
  XOR2_X1 U401 ( .A(G162GAT), .B(KEYINPUT74), .Z(n385) );
  XNOR2_X1 U402 ( .A(n377), .B(n385), .ZN(n340) );
  XOR2_X1 U403 ( .A(KEYINPUT21), .B(G211GAT), .Z(n339) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(G218GAT), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n419) );
  XOR2_X1 U406 ( .A(n344), .B(n343), .Z(n468) );
  XOR2_X1 U407 ( .A(KEYINPUT47), .B(KEYINPUT115), .Z(n404) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(G211GAT), .Z(n346) );
  XNOR2_X1 U409 ( .A(G183GAT), .B(KEYINPUT12), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U411 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U412 ( .A(KEYINPUT79), .B(KEYINPUT77), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n364) );
  XOR2_X1 U415 ( .A(G155GAT), .B(G127GAT), .Z(n352) );
  XNOR2_X1 U416 ( .A(G22GAT), .B(G8GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U418 ( .A(G64GAT), .B(G78GAT), .Z(n354) );
  XNOR2_X1 U419 ( .A(G15GAT), .B(G71GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U421 ( .A(n356), .B(n355), .Z(n362) );
  XOR2_X1 U422 ( .A(G1GAT), .B(KEYINPUT69), .Z(n368) );
  XOR2_X1 U423 ( .A(n357), .B(KEYINPUT78), .Z(n359) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n368), .B(n360), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n570) );
  XOR2_X1 U429 ( .A(G29GAT), .B(G50GAT), .Z(n366) );
  XNOR2_X1 U430 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n391) );
  XNOR2_X1 U432 ( .A(n391), .B(KEYINPUT30), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n367), .B(G197GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n368), .B(KEYINPUT68), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n369), .B(KEYINPUT29), .ZN(n370) );
  XOR2_X1 U436 ( .A(n371), .B(n370), .Z(n375) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(G36GAT), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n372), .B(G8GAT), .ZN(n412) );
  XNOR2_X1 U439 ( .A(n412), .B(n373), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U441 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U442 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n576) );
  NOR2_X1 U444 ( .A1(n576), .A2(n558), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n380), .B(KEYINPUT46), .ZN(n381) );
  NOR2_X1 U446 ( .A1(n570), .A2(n381), .ZN(n402) );
  XOR2_X1 U447 ( .A(G106GAT), .B(KEYINPUT10), .Z(n383) );
  XNOR2_X1 U448 ( .A(G99GAT), .B(KEYINPUT76), .ZN(n382) );
  XOR2_X1 U449 ( .A(n383), .B(n382), .Z(n401) );
  XOR2_X1 U450 ( .A(G218GAT), .B(n384), .Z(n387) );
  XNOR2_X1 U451 ( .A(G43GAT), .B(n385), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n393) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n389) );
  XOR2_X1 U454 ( .A(n393), .B(n392), .Z(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT66), .B(KEYINPUT75), .Z(n395) );
  XNOR2_X1 U456 ( .A(G36GAT), .B(KEYINPUT9), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n566) );
  NAND2_X1 U461 ( .A1(n402), .A2(n566), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n409) );
  XOR2_X1 U463 ( .A(n576), .B(KEYINPUT70), .Z(n568) );
  INV_X1 U464 ( .A(n570), .ZN(n584) );
  XNOR2_X1 U465 ( .A(n566), .B(KEYINPUT36), .ZN(n587) );
  NOR2_X1 U466 ( .A1(n584), .A2(n587), .ZN(n405) );
  NOR2_X1 U467 ( .A1(n481), .A2(n297), .ZN(n406) );
  XOR2_X1 U468 ( .A(KEYINPUT116), .B(n406), .Z(n407) );
  NOR2_X1 U469 ( .A1(n568), .A2(n407), .ZN(n408) );
  XNOR2_X1 U470 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n553) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(n412), .Z(n414) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U475 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n416) );
  XNOR2_X1 U476 ( .A(G190GAT), .B(G92GAT), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U478 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n483) );
  NOR2_X1 U482 ( .A1(n553), .A2(n483), .ZN(n426) );
  XNOR2_X1 U483 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n448) );
  XOR2_X1 U485 ( .A(KEYINPUT90), .B(KEYINPUT76), .Z(n428) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(G113GAT), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U488 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n430) );
  XNOR2_X1 U489 ( .A(G120GAT), .B(KEYINPUT6), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U491 ( .A(n432), .B(n431), .Z(n438) );
  XOR2_X1 U492 ( .A(G162GAT), .B(n433), .Z(n435) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(G85GAT), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U495 ( .A(G134GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n447) );
  XOR2_X1 U497 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n440) );
  XNOR2_X1 U498 ( .A(G1GAT), .B(G57GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n445) );
  XOR2_X1 U500 ( .A(n441), .B(G148GAT), .Z(n443) );
  NAND2_X1 U501 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U503 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n526) );
  NAND2_X1 U505 ( .A1(n448), .A2(n526), .ZN(n449) );
  XOR2_X1 U506 ( .A(n449), .B(KEYINPUT65), .Z(n573) );
  NOR2_X1 U507 ( .A1(n468), .A2(n573), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NAND2_X1 U509 ( .A1(n540), .A2(n571), .ZN(n455) );
  XOR2_X1 U510 ( .A(G176GAT), .B(KEYINPUT125), .Z(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  INV_X1 U514 ( .A(n566), .ZN(n547) );
  NAND2_X1 U515 ( .A1(n571), .A2(n547), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n457) );
  INV_X1 U517 ( .A(G190GAT), .ZN(n456) );
  NOR2_X1 U518 ( .A1(n536), .A2(n483), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n468), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT25), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n463) );
  NAND2_X1 U522 ( .A1(n468), .A2(n536), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n574) );
  XOR2_X1 U524 ( .A(KEYINPUT27), .B(n483), .Z(n470) );
  NAND2_X1 U525 ( .A1(n574), .A2(n470), .ZN(n552) );
  NAND2_X1 U526 ( .A1(n464), .A2(n552), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n465), .A2(n526), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT95), .ZN(n474) );
  INV_X1 U529 ( .A(n526), .ZN(n555) );
  INV_X1 U530 ( .A(KEYINPUT67), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n535) );
  XNOR2_X1 U533 ( .A(n536), .B(KEYINPUT85), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n535), .A2(n472), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n475), .B(KEYINPUT96), .ZN(n489) );
  NOR2_X1 U537 ( .A1(n570), .A2(n489), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n476), .B(KEYINPUT101), .ZN(n477) );
  NOR2_X1 U539 ( .A1(n587), .A2(n477), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n478) );
  INV_X1 U541 ( .A(n481), .ZN(n580) );
  NAND2_X1 U542 ( .A1(n568), .A2(n580), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n525), .A2(n491), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT38), .B(n482), .Z(n509) );
  NOR2_X1 U545 ( .A1(n509), .A2(n483), .ZN(n486) );
  NOR2_X1 U546 ( .A1(n547), .A2(n584), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NOR2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT97), .B(n490), .ZN(n512) );
  OR2_X1 U550 ( .A1(n491), .A2(n512), .ZN(n500) );
  NOR2_X1 U551 ( .A1(n526), .A2(n500), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT98), .B(KEYINPUT34), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U554 ( .A(G1GAT), .B(n494), .Z(G1324GAT) );
  NOR2_X1 U555 ( .A1(n483), .A2(n500), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U558 ( .A1(n536), .A2(n500), .ZN(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n532), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(G22GAT), .B(n501), .Z(G1327GAT) );
  NOR2_X1 U564 ( .A1(n526), .A2(n509), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n503) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XNOR2_X1 U569 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n507) );
  NOR2_X1 U570 ( .A1(n536), .A2(n509), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n532), .A2(n509), .ZN(n510) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  NAND2_X1 U575 ( .A1(n540), .A2(n576), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(KEYINPUT110), .ZN(n524) );
  NOR2_X1 U577 ( .A1(n512), .A2(n524), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT111), .ZN(n521) );
  NOR2_X1 U579 ( .A1(n526), .A2(n521), .ZN(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U582 ( .A(G57GAT), .B(n516), .Z(G1332GAT) );
  NOR2_X1 U583 ( .A1(n483), .A2(n521), .ZN(n517) );
  XOR2_X1 U584 ( .A(KEYINPUT112), .B(n517), .Z(n518) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n536), .A2(n521), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G71GAT), .B(KEYINPUT113), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1334GAT) );
  NOR2_X1 U589 ( .A1(n532), .A2(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  OR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U593 ( .A1(n526), .A2(n531), .ZN(n527) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n483), .A2(n531), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(n528), .Z(n529) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n536), .A2(n531), .ZN(n530) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT117), .Z(n539) );
  OR2_X1 U604 ( .A1(n536), .A2(n553), .ZN(n537) );
  NOR2_X1 U605 ( .A1(n535), .A2(n537), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n548), .A2(n568), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U609 ( .A1(n548), .A2(n540), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n544) );
  NAND2_X1 U613 ( .A1(n548), .A2(n570), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(n556), .Z(n565) );
  NOR2_X1 U623 ( .A1(n576), .A2(n565), .ZN(n557) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n557), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n565), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n560) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT122), .B(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n584), .A2(n565), .ZN(n564) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n571), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U639 ( .A(n573), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n576), .A2(n586), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n586), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

