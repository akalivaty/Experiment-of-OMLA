//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(new_n448), .B2(new_n456), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n467), .A3(G137), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  XNOR2_X1  g051(.A(KEYINPUT67), .B(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n467), .A2(new_n472), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G124), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n487), .A3(G2104), .ZN(new_n488));
  AND2_X1   g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G138), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n494), .B2(new_n477), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n466), .A2(new_n467), .A3(new_n496), .A4(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .A3(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g083(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  XOR2_X1   g087(.A(new_n512), .B(KEYINPUT69), .Z(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n501), .A2(new_n503), .B1(KEYINPUT6), .B2(new_n500), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(G50), .A3(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n510), .A2(new_n514), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  XNOR2_X1  g093(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n519));
  AND3_X1   g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(new_n522), .B1(new_n508), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n509), .A2(G89), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(G543), .B1(new_n515), .B2(KEYINPUT70), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n504), .A2(KEYINPUT70), .A3(new_n505), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n529), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n506), .A2(new_n507), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(G90), .B1(new_n537), .B2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  XNOR2_X1  g115(.A(KEYINPUT72), .B(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n509), .A2(G81), .B1(new_n545), .B2(G651), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  XNOR2_X1  g127(.A(KEYINPUT73), .B(G65), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(new_n508), .B1(G78), .B2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT74), .B1(new_n555), .B2(new_n500), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(new_n535), .B2(new_n553), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(new_n559), .A3(G651), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n556), .A2(new_n560), .B1(G91), .B2(new_n509), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n529), .B2(G53), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  NOR4_X1   g139(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT9), .A4(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(G299));
  OAI21_X1  g141(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n504), .A2(new_n505), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(G543), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n571), .B1(new_n576), .B2(new_n577), .ZN(G288));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n506), .B2(new_n507), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n504), .A2(G86), .A3(new_n508), .A4(new_n505), .ZN(new_n584));
  AND2_X1   g159(.A1(G48), .A2(G543), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n504), .A2(new_n505), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n529), .A2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n535), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n509), .A2(G85), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n509), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n574), .A2(G54), .A3(G543), .A4(new_n575), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI211_X1 g175(.A(KEYINPUT75), .B(new_n599), .C1(new_n535), .C2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n600), .B1(new_n506), .B2(new_n507), .ZN(new_n603));
  INV_X1    g178(.A(new_n599), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n601), .A2(new_n605), .A3(G651), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n597), .A2(new_n598), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n598), .B1(new_n597), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n596), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT77), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G171), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT78), .Z(G284));
  INV_X1    g190(.A(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G299), .A2(new_n611), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n611), .B2(G168), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n610), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n467), .A2(new_n473), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n479), .A2(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n480), .A2(G135), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  INV_X1    g237(.A(new_n656), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n658), .A3(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n657), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n679), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n683));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n675), .A2(new_n684), .A3(new_n678), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n684), .B1(new_n675), .B2(new_n678), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n675), .A2(new_n678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(KEYINPUT81), .ZN(new_n690));
  INV_X1    g265(.A(new_n683), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n682), .A2(new_n688), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n682), .A2(new_n688), .A3(KEYINPUT82), .A4(new_n692), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n672), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(new_n697), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G1981), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n703), .A2(G1986), .A3(new_n698), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT83), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n701), .B2(new_n704), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n671), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n699), .A2(new_n700), .A3(new_n672), .ZN(new_n711));
  AOI21_X1  g286(.A(G1986), .B1(new_n703), .B2(new_n698), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(new_n670), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n715), .ZN(G229));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G26), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n479), .A2(G128), .B1(new_n480), .B2(G140), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT88), .B(G2067), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2072), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n719), .A2(G33), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(new_n466), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G139), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n729), .B1(new_n736), .B2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n727), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n483), .A2(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n719), .A2(G35), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n742), .A2(new_n743), .A3(G2090), .ZN(new_n744));
  AND2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n719), .B1(KEYINPUT24), .B2(G34), .ZN(new_n746));
  OAI22_X1  g321(.A1(G160), .A2(new_n719), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(G2084), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(G2084), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n635), .A2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n751), .A2(new_n719), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND4_X1   g329(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(G2090), .B1(new_n742), .B2(new_n743), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n738), .A2(new_n744), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n737), .A2(new_n728), .B1(G2078), .B2(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G19), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n547), .B2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(G1341), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n478), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n473), .A2(G105), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n467), .A2(new_n472), .ZN(new_n772));
  INV_X1    g347(.A(G141), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR3_X1    g349(.A1(new_n770), .A2(new_n774), .A3(KEYINPUT89), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT89), .B1(new_n770), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n775), .A2(KEYINPUT90), .A3(new_n776), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n719), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT91), .ZN(new_n784));
  NOR2_X1   g359(.A1(G29), .A2(G32), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n782), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n782), .B2(new_n786), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n757), .A2(new_n765), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G16), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n610), .B2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1348), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT93), .B(KEYINPUT23), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n790), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NOR2_X1   g373(.A1(G5), .A2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G171), .B2(G16), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1961), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n764), .A2(G1341), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n790), .A2(G21), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G286), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(G1966), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n800), .A2(G1961), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n801), .A2(new_n802), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n805), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT92), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n789), .A2(new_n793), .A3(new_n798), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n792), .A2(G1348), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n717), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n757), .A2(new_n765), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n787), .A2(new_n788), .ZN(new_n816));
  AND4_X1   g391(.A1(new_n798), .A2(new_n815), .A3(new_n816), .A4(new_n811), .ZN(new_n817));
  INV_X1    g392(.A(new_n813), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n817), .A2(KEYINPUT94), .A3(new_n818), .A4(new_n793), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n790), .A2(G22), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G166), .B2(new_n790), .ZN(new_n823));
  INV_X1    g398(.A(G1971), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n790), .A2(G23), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n570), .B1(new_n529), .B2(G49), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n790), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT33), .B(G1976), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT86), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  MUX2_X1   g407(.A(G6), .B(G305), .S(G16), .Z(new_n833));
  XOR2_X1   g408(.A(KEYINPUT32), .B(G1981), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n825), .A2(new_n831), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT34), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n790), .A2(G24), .ZN(new_n838));
  INV_X1    g413(.A(G290), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n790), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n672), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT85), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n719), .A2(G25), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT84), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n479), .A2(G119), .B1(new_n480), .B2(G131), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n845), .B1(new_n850), .B2(new_n719), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT35), .B(G1991), .Z(new_n852));
  XOR2_X1   g427(.A(new_n851), .B(new_n852), .Z(new_n853));
  NOR2_X1   g428(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n837), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n820), .A2(new_n821), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n821), .B1(new_n820), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(G311));
  NAND2_X1  g434(.A1(new_n820), .A2(new_n856), .ZN(G150));
  NAND2_X1  g435(.A1(new_n610), .A2(G559), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n542), .B2(new_n546), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n509), .A2(G93), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n500), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT97), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n866), .A2(new_n869), .A3(new_n500), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT98), .B(G55), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n576), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n542), .A2(new_n862), .A3(new_n546), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n864), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n865), .B1(new_n576), .B2(new_n872), .C1(new_n868), .C2(new_n870), .ZN(new_n877));
  INV_X1    g452(.A(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n863), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n861), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g459(.A(G860), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n877), .A2(G860), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G145));
  NAND2_X1  g464(.A1(new_n849), .A2(new_n627), .ZN(new_n890));
  INV_X1    g465(.A(new_n627), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n847), .A2(new_n891), .A3(new_n848), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n480), .A2(G142), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT101), .Z(new_n895));
  NOR2_X1   g470(.A1(new_n466), .A2(G118), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  INV_X1    g472(.A(G130), .ZN(new_n898));
  OAI22_X1  g473(.A1(new_n896), .A2(new_n897), .B1(new_n478), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n890), .A3(new_n892), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n495), .A2(new_n497), .ZN(new_n908));
  INV_X1    g483(.A(new_n493), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n736), .B1(new_n779), .B2(new_n780), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n777), .A2(new_n736), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n724), .B(KEYINPUT100), .ZN(new_n915));
  INV_X1    g490(.A(new_n736), .ZN(new_n916));
  INV_X1    g491(.A(new_n780), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT90), .B1(new_n775), .B2(new_n776), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(G164), .A3(new_n912), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n915), .B1(new_n914), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n914), .A2(new_n920), .ZN(new_n924));
  INV_X1    g499(.A(new_n915), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n914), .A2(new_n920), .A3(new_n915), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n906), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n635), .B(G160), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(new_n483), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n923), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n923), .B2(new_n928), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n931), .A2(new_n932), .A3(G37), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT40), .Z(G395));
  OAI211_X1 g509(.A(new_n609), .B(new_n561), .C1(new_n563), .C2(new_n565), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n594), .B(KEYINPUT10), .ZN(new_n937));
  INV_X1    g512(.A(new_n608), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n597), .A2(new_n598), .A3(new_n606), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G299), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(KEYINPUT103), .A3(G299), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n935), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(KEYINPUT41), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n622), .B(new_n880), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n950), .B2(new_n947), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n827), .B(G305), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g529(.A1(G303), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT104), .A4(new_n516), .ZN(new_n956));
  NAND3_X1  g531(.A1(G290), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G290), .B1(new_n955), .B2(new_n956), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(G288), .B(G305), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(new_n956), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n839), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n963), .A3(new_n957), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n964), .A3(KEYINPUT105), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n952), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n952), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(G868), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G868), .B2(new_n874), .ZN(G295));
  OAI21_X1  g546(.A(new_n970), .B1(G868), .B2(new_n874), .ZN(G331));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n960), .A2(new_n964), .ZN(new_n974));
  NOR2_X1   g549(.A1(G286), .A2(G301), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n530), .A2(new_n526), .B1(new_n533), .B2(new_n538), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n977), .A2(new_n876), .A3(new_n879), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n876), .B2(new_n879), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n947), .A2(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(new_n942), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n947), .A2(new_n978), .A3(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G37), .ZN(new_n985));
  INV_X1    g560(.A(new_n947), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n980), .B2(new_n936), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n974), .B(KEYINPUT107), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n935), .A2(new_n941), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT41), .B(new_n989), .C1(new_n978), .C2(new_n979), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n984), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n973), .B1(new_n992), .B2(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n980), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n988), .B(new_n994), .C1(new_n948), .C2(new_n980), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n984), .A2(new_n995), .A3(new_n985), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n993), .B1(KEYINPUT43), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n984), .A2(new_n991), .A3(new_n999), .A4(new_n985), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT108), .B1(new_n1001), .B2(new_n973), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n1003), .B(KEYINPUT44), .C1(new_n998), .C2(new_n1000), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(G397));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(G164), .B2(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n468), .A2(new_n469), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n477), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(G40), .A3(new_n474), .A4(new_n471), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n839), .A2(new_n672), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n917), .B2(new_n918), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n850), .A2(new_n852), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n724), .A2(G2067), .ZN(new_n1017));
  INV_X1    g592(.A(G2067), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n722), .A2(new_n1018), .A3(new_n723), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(G1996), .B2(new_n777), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n850), .A2(new_n852), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1015), .A2(new_n1016), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1011), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1013), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1025), .B2(G1996), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1011), .A2(KEYINPUT46), .A3(new_n1014), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1011), .B1(new_n1020), .B2(new_n777), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1019), .B1(new_n1033), .B2(new_n1022), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1011), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1026), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n910), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1010), .B1(new_n1038), .B2(new_n1006), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT56), .B(G2072), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n910), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT109), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G164), .A2(G1384), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT45), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1039), .B(new_n1040), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n561), .B(new_n1048), .C1(new_n563), .C2(new_n565), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n910), .A2(new_n1050), .A3(new_n1037), .ZN(new_n1051));
  INV_X1    g626(.A(G40), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n470), .A2(new_n475), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1956), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1046), .A2(new_n1057), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1059));
  INV_X1    g634(.A(G1348), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1038), .A2(new_n1010), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1055), .A2(new_n1060), .B1(new_n1061), .B2(new_n1018), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n609), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1058), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1046), .A2(new_n1057), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(KEYINPUT120), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1058), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(KEYINPUT120), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(G1341), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1007), .A2(new_n1053), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1041), .A2(KEYINPUT109), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1044), .A2(new_n1043), .A3(KEYINPUT45), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1085), .B2(new_n1014), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n542), .A2(new_n546), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT59), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1014), .B(new_n1039), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1080), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n547), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1075), .A2(KEYINPUT61), .A3(new_n1058), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1061), .A2(new_n1018), .ZN(new_n1096));
  AND4_X1   g671(.A1(KEYINPUT60), .A2(new_n1095), .A3(new_n609), .A4(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n609), .B1(new_n1062), .B2(KEYINPUT60), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1093), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1066), .B(new_n1067), .C1(new_n1076), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G2078), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1085), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(KEYINPUT122), .A3(new_n1105), .ZN(new_n1109));
  INV_X1    g684(.A(G1961), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1055), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n475), .B(KEYINPUT123), .Z(new_n1112));
  NAND3_X1  g687(.A1(new_n1103), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1112), .A2(new_n470), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1114), .B(new_n1007), .C1(new_n1045), .C2(new_n1042), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1106), .A2(new_n1107), .B1(new_n1110), .B2(new_n1055), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1082), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1120), .A2(new_n1041), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1007), .A2(KEYINPUT117), .A3(new_n1053), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1103), .A4(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1041), .A3(new_n1123), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n1125), .B2(G2078), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(KEYINPUT53), .A3(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1118), .A2(new_n1127), .A3(G301), .A4(new_n1109), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1117), .A2(new_n1128), .A3(KEYINPUT54), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n571), .B(G1976), .C1(new_n576), .C2(new_n577), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1077), .A3(G8), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n827), .B2(G1976), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT111), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1976), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT52), .B1(G288), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT111), .ZN(new_n1137));
  INV_X1    g712(.A(G8), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .A4(new_n1130), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n583), .A2(new_n584), .A3(new_n696), .A4(new_n586), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT112), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1143), .B(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n508), .A2(G61), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n500), .B1(new_n1146), .B2(new_n581), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n584), .A2(new_n586), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(KEYINPUT113), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT113), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n584), .A2(new_n1150), .A3(new_n586), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n696), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1142), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1143), .B(KEYINPUT112), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1148), .A2(KEYINPUT113), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n583), .A3(new_n1151), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G1981), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1157), .A3(KEYINPUT49), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1158), .A3(new_n1139), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1131), .A2(KEYINPUT52), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1141), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G303), .A2(G8), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT55), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1085), .A2(G1971), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT110), .B(G2090), .Z(new_n1166));
  NOR2_X1   g741(.A1(new_n1055), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1164), .B(G8), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1039), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1169), .B2(new_n824), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1163), .B1(new_n1170), .B2(new_n1138), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1161), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1055), .A2(G2084), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1125), .B2(new_n805), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1138), .B1(new_n1174), .B2(G168), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT51), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT51), .B1(new_n1174), .B2(G168), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1175), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1172), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1116), .A2(G301), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1118), .A2(new_n1127), .A3(G171), .A4(new_n1109), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1102), .A2(new_n1129), .A3(new_n1180), .A4(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1170), .A2(new_n1138), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1134), .A2(new_n1140), .B1(KEYINPUT52), .B2(new_n1131), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1186), .A2(new_n1159), .A3(new_n1187), .A4(new_n1164), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1139), .B(KEYINPUT114), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G288), .A2(G1976), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1145), .B1(new_n1159), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT115), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g768(.A(KEYINPUT115), .B(new_n1145), .C1(new_n1159), .C2(new_n1190), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(KEYINPUT116), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT116), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1188), .B(new_n1197), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n1199));
  NAND2_X1  g774(.A1(G168), .A2(G8), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1174), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1199), .B1(new_n1172), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1171), .A2(new_n1168), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1204), .A2(KEYINPUT63), .A3(new_n1161), .A4(new_n1201), .ZN(new_n1205));
  AOI22_X1  g780(.A1(new_n1196), .A2(new_n1198), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1185), .A2(KEYINPUT124), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT124), .B1(new_n1185), .B2(new_n1206), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1177), .A2(new_n1209), .A3(new_n1179), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1172), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1118), .A2(new_n1127), .A3(new_n1109), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1210), .A2(new_n1211), .A3(G171), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1214), .B1(new_n1215), .B2(KEYINPUT62), .ZN(new_n1216));
  AOI211_X1 g791(.A(KEYINPUT125), .B(new_n1209), .C1(new_n1177), .C2(new_n1179), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1213), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1207), .A2(new_n1208), .A3(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(G290), .B(new_n672), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1025), .B1(new_n1024), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1036), .B1(new_n1219), .B2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g797(.A1(new_n462), .A2(G227), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n653), .A2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g799(.A(new_n1225), .B(KEYINPUT126), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n710), .A2(new_n715), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g801(.A1(new_n933), .A2(new_n1227), .ZN(new_n1228));
  AND3_X1   g802(.A1(new_n1228), .A2(new_n1001), .A3(KEYINPUT127), .ZN(new_n1229));
  AOI21_X1  g803(.A(KEYINPUT127), .B1(new_n1228), .B2(new_n1001), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1229), .A2(new_n1230), .ZN(G308));
  NAND2_X1  g805(.A1(new_n1228), .A2(new_n1001), .ZN(G225));
endmodule


