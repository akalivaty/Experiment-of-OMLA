//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT23), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT24), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n209), .A2(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(KEYINPUT24), .B2(new_n204), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n203), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT66), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT27), .B(G183gat), .Z(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n225));
  AOI21_X1  g024(.A(G190gat), .B1(new_n225), .B2(KEYINPUT65), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT28), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n222), .A2(new_n228), .A3(G190gat), .ZN(new_n229));
  OAI221_X1 g028(.A(new_n204), .B1(new_n216), .B2(new_n221), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n231), .A2(G226gat), .A3(G233gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n231), .A2(new_n233), .B1(G226gat), .B2(G233gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT70), .B(G197gat), .ZN(new_n236));
  INV_X1    g035(.A(G204gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  INV_X1    g038(.A(G211gat), .ZN(new_n240));
  INV_X1    g039(.A(G218gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n238), .A2(new_n239), .B1(KEYINPUT22), .B2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G211gat), .B(G218gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n232), .A2(new_n234), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G8gat), .B(G36gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT71), .ZN(new_n251));
  XNOR2_X1  g050(.A(G64gat), .B(G92gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT30), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  INV_X1    g058(.A(new_n253), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n246), .B2(new_n248), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G113gat), .B(G120gat), .Z(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271));
  XOR2_X1   g070(.A(G141gat), .B(G148gat), .Z(new_n272));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G162gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(G155gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G162gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT73), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n272), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(G162gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n273), .B1(new_n285), .B2(G155gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n280), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OR3_X1    g086(.A1(new_n270), .A2(new_n271), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n271), .B1(new_n270), .B2(new_n287), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n270), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT5), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n270), .B(new_n287), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n295), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n298), .A2(new_n299), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G1gat), .B(G29gat), .Z(new_n304));
  XNOR2_X1  g103(.A(G57gat), .B(G85gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n311), .B(KEYINPUT39), .C1(new_n295), .C2(new_n301), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(new_n308), .C1(KEYINPUT39), .C2(new_n311), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT40), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n262), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n303), .A2(new_n317), .A3(new_n308), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n303), .B2(new_n308), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n310), .B(new_n316), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  OR3_X1    g119(.A1(new_n246), .A2(KEYINPUT37), .A3(new_n248), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT37), .B1(new_n246), .B2(new_n248), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n260), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(KEYINPUT38), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(KEYINPUT38), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n324), .A2(new_n254), .A3(new_n325), .ZN(new_n326));
  OR3_X1    g125(.A1(new_n303), .A2(new_n308), .A3(new_n316), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n315), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n245), .A2(new_n233), .A3(new_n287), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n287), .A2(new_n291), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT82), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n292), .A2(new_n233), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n247), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n334), .A2(KEYINPUT82), .ZN(new_n339));
  INV_X1    g138(.A(G228gat), .ZN(new_n340));
  INV_X1    g139(.A(G233gat), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n290), .A2(new_n340), .A3(new_n341), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n332), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G22gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  INV_X1    g146(.A(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G22gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n351), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n350), .B1(new_n346), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n331), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n330), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n231), .B1(KEYINPUT68), .B2(new_n270), .ZN(new_n363));
  INV_X1    g162(.A(new_n270), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n231), .A2(new_n365), .A3(new_n364), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n367), .A2(G227gat), .A3(G233gat), .A4(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n368), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT34), .ZN(new_n373));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  OR3_X1    g175(.A1(new_n371), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n371), .A2(new_n375), .A3(new_n376), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n385), .A2(KEYINPUT69), .A3(KEYINPUT36), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT36), .B1(new_n385), .B2(KEYINPUT69), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n329), .A2(new_n359), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT35), .ZN(new_n390));
  INV_X1    g189(.A(new_n262), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n356), .B2(new_n358), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n320), .A2(new_n327), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n359), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n388), .A2(new_n396), .B1(KEYINPUT35), .B2(new_n392), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n309), .B(KEYINPUT80), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n327), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n391), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n389), .B(new_n395), .C1(new_n397), .C2(new_n401), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n348), .A2(G43gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n348), .A2(G43gat), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n403), .A2(KEYINPUT15), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT84), .B(G43gat), .Z(new_n407));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n348), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT84), .B(G43gat), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT85), .B1(new_n410), .B2(G50gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n403), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT15), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT14), .B(G29gat), .Z(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(G36gat), .ZN(new_n416));
  INV_X1    g215(.A(G29gat), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n417), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n406), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G8gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G15gat), .B(G22gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(G1gat), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(KEYINPUT87), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(G1gat), .B2(new_n422), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n405), .B1(new_n416), .B2(new_n418), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n420), .A2(new_n431), .A3(KEYINPUT17), .A4(new_n428), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n419), .B1(new_n412), .B2(new_n413), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n431), .B(new_n428), .C1(new_n433), .C2(new_n405), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n427), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G229gat), .A2(G233gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(KEYINPUT18), .A3(new_n440), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n440), .B(KEYINPUT13), .Z(new_n445));
  AOI21_X1  g244(.A(new_n427), .B1(new_n420), .B2(new_n428), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n430), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT88), .B(new_n445), .C1(new_n430), .C2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n443), .A2(new_n444), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(G169gat), .B(G197gat), .Z(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n451), .A4(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n402), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT89), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n402), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n400), .ZN(new_n468));
  INV_X1    g267(.A(G92gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G92gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT94), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(G99gat), .A3(G106gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT8), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G99gat), .B(G106gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(new_n479), .A3(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n437), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(G190gat), .B(G218gat), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT41), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n420), .A2(new_n428), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n486), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n485), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n432), .B2(new_n436), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n487), .B1(new_n497), .B2(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n490), .A2(KEYINPUT41), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(KEYINPUT93), .Z(new_n501));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n495), .A2(new_n503), .A3(new_n498), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G57gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G57gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(G64gat), .ZN(new_n512));
  INV_X1    g311(.A(G64gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G57gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G71gat), .ZN(new_n516));
  INV_X1    g315(.A(G78gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT9), .ZN(new_n518));
  NAND2_X1  g317(.A1(G71gat), .A2(G78gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n508), .A2(G64gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT9), .ZN(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G78gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n515), .A2(new_n520), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n427), .B1(KEYINPUT21), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(KEYINPUT21), .ZN(new_n528));
  XNOR2_X1  g327(.A(G127gat), .B(G155gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n527), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT91), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT92), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n531), .B(new_n538), .Z(new_n539));
  NOR2_X1   g338(.A1(new_n507), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G230gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n341), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n483), .A3(new_n484), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n474), .A2(new_n481), .A3(new_n479), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n481), .B1(new_n474), .B2(new_n479), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n512), .A2(new_n514), .B1(new_n519), .B2(new_n518), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n524), .B1(KEYINPUT9), .B2(new_n522), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n526), .A2(new_n483), .A3(KEYINPUT95), .A4(new_n484), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT10), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554));
  INV_X1    g353(.A(new_n544), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n553), .A2(new_n554), .B1(KEYINPUT10), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n552), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT10), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT96), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n543), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n543), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n561), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n541), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n467), .A2(new_n468), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G1gat), .ZN(G1324gat));
  INV_X1    g374(.A(new_n573), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(new_n464), .B2(new_n466), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n262), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT42), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT97), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT16), .B(G8gat), .Z(new_n581));
  MUX2_X1   g380(.A(KEYINPUT97), .B(new_n580), .S(new_n581), .Z(new_n582));
  NOR2_X1   g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n578), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n579), .B1(new_n584), .B2(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(G8gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(G1325gat));
  INV_X1    g386(.A(G15gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n385), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n577), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n386), .A2(new_n387), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n577), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n592), .B2(new_n588), .ZN(G1326gat));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n396), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT43), .B(G22gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(G1327gat));
  INV_X1    g395(.A(new_n572), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n539), .ZN(new_n598));
  INV_X1    g397(.A(new_n507), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n467), .A2(new_n417), .A3(new_n468), .A4(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT98), .B(KEYINPUT45), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n402), .A2(new_n604), .A3(new_n507), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT44), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n402), .A2(new_n604), .A3(KEYINPUT44), .A4(new_n507), .ZN(new_n608));
  INV_X1    g407(.A(new_n462), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n598), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n607), .A2(new_n468), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n417), .B1(new_n611), .B2(KEYINPUT100), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(KEYINPUT100), .B2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n613), .ZN(G1328gat));
  INV_X1    g413(.A(new_n600), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n464), .B2(new_n466), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n391), .A2(G36gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OR3_X1    g418(.A1(new_n617), .A2(KEYINPUT46), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT46), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  INV_X1    g420(.A(G36gat), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n607), .A2(new_n608), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n623), .A2(new_n262), .A3(new_n610), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n624), .ZN(G1329gat));
  NAND4_X1  g424(.A1(new_n607), .A2(new_n591), .A3(new_n608), .A4(new_n610), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n407), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n589), .A2(new_n410), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n617), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT47), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n627), .B(KEYINPUT47), .C1(new_n617), .C2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(G1330gat));
  INV_X1    g432(.A(KEYINPUT48), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n359), .A2(G50gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT101), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n616), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n607), .A2(new_n396), .A3(new_n608), .A4(new_n610), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(G50gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n638), .A2(G50gat), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n616), .A2(new_n636), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n634), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(G1331gat));
  NOR3_X1   g445(.A1(new_n541), .A2(new_n462), .A3(new_n597), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n402), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n468), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n509), .A2(new_n511), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1332gat));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n402), .A2(KEYINPUT103), .A3(new_n647), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n262), .B(KEYINPUT104), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT105), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n654), .A2(new_n660), .A3(new_n655), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1333gat));
  NAND2_X1  g463(.A1(new_n654), .A2(new_n655), .ZN(new_n665));
  OAI21_X1  g464(.A(G71gat), .B1(new_n665), .B2(new_n388), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n516), .A3(new_n589), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT50), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1334gat));
  NOR2_X1   g469(.A1(new_n665), .A2(new_n359), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n517), .ZN(G1335gat));
  INV_X1    g471(.A(new_n539), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n462), .A2(new_n673), .A3(new_n597), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n623), .A2(new_n468), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G85gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n462), .A2(new_n673), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n402), .A2(new_n507), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT51), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT51), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n402), .A2(new_n680), .A3(new_n507), .A4(new_n677), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n572), .A3(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n400), .A2(G85gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(G1336gat));
  INV_X1    g483(.A(new_n682), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n656), .A2(G92gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT52), .ZN(new_n688));
  INV_X1    g487(.A(new_n656), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n607), .A2(new_n608), .A3(new_n689), .A4(new_n674), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G92gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n607), .A2(new_n262), .A3(new_n608), .A4(new_n674), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n685), .A2(new_n686), .B1(new_n693), .B2(G92gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n688), .B2(new_n694), .ZN(G1337gat));
  NAND3_X1  g494(.A1(new_n623), .A2(new_n591), .A3(new_n674), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G99gat), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n385), .A2(G99gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n682), .B2(new_n698), .ZN(G1338gat));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n359), .A2(G106gat), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n682), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT53), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n607), .A2(new_n396), .A3(new_n608), .A4(new_n674), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G106gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT53), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1339gat));
  INV_X1    g510(.A(KEYINPUT55), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT54), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n556), .A2(new_n560), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n563), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n556), .A2(new_n560), .A3(new_n543), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n557), .A2(new_n554), .A3(new_n558), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n555), .A2(KEYINPUT10), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n553), .A2(new_n554), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n713), .B(new_n563), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(new_n723), .A3(new_n570), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n722), .B2(new_n570), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n717), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n717), .B(new_n728), .C1(new_n724), .C2(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n569), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n724), .B2(new_n725), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(new_n712), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n430), .A2(new_n446), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n439), .A2(new_n440), .B1(new_n735), .B2(new_n445), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n457), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n507), .A2(new_n461), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n730), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n730), .A2(new_n741), .A3(new_n734), .A4(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n461), .A2(new_n572), .A3(new_n737), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT110), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n462), .A3(new_n734), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n507), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n539), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n573), .A2(new_n609), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n396), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n750), .A2(new_n589), .A3(new_n468), .A4(new_n656), .ZN(new_n751));
  INV_X1    g550(.A(G113gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n609), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n400), .B1(new_n748), .B2(new_n749), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n392), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n656), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n462), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n757), .B2(new_n752), .ZN(G1340gat));
  INV_X1    g557(.A(G120gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(new_n759), .A3(new_n572), .ZN(new_n760));
  OAI21_X1  g559(.A(G120gat), .B1(new_n751), .B2(new_n597), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT111), .Z(G1341gat));
  INV_X1    g562(.A(G127gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n756), .A2(new_n764), .A3(new_n673), .ZN(new_n765));
  OAI21_X1  g564(.A(G127gat), .B1(new_n751), .B2(new_n539), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1342gat));
  INV_X1    g566(.A(G134gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n262), .A2(new_n599), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n755), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n770), .A2(KEYINPUT56), .ZN(new_n771));
  OAI21_X1  g570(.A(G134gat), .B1(new_n751), .B2(new_n599), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(KEYINPUT56), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(G1343gat));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n754), .A2(new_n396), .A3(new_n388), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n609), .A2(G141gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT115), .Z(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n656), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n689), .A2(new_n591), .A3(new_n400), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n396), .A2(KEYINPUT57), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n731), .B1(new_n733), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n729), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n722), .A2(new_n570), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT107), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n722), .A2(new_n723), .A3(new_n570), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n728), .B1(new_n789), .B2(new_n717), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT113), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n730), .A2(new_n793), .A3(new_n784), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n462), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n507), .B1(new_n795), .B2(new_n744), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n539), .B1(new_n796), .B2(new_n743), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n782), .B1(new_n797), .B2(new_n749), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n748), .A2(new_n749), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT57), .B1(new_n799), .B2(new_n396), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n462), .B(new_n781), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G141gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n780), .B1(new_n802), .B2(KEYINPUT114), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n804), .A3(G141gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n776), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n780), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n775), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n801), .A2(new_n804), .A3(G141gat), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n804), .B1(new_n801), .B2(G141gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(new_n780), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT117), .B(new_n809), .C1(new_n814), .C2(new_n776), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(G1344gat));
  AND2_X1   g615(.A1(new_n777), .A2(new_n656), .ZN(new_n817));
  INV_X1    g616(.A(G148gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n572), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n799), .A2(KEYINPUT57), .A3(new_n396), .ZN(new_n821));
  INV_X1    g620(.A(new_n739), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n539), .B1(new_n796), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n359), .B1(new_n823), .B2(new_n749), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n821), .B1(new_n824), .B2(KEYINPUT57), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n825), .A2(new_n572), .A3(new_n781), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n818), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n820), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n781), .B1(new_n798), .B2(new_n800), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(new_n597), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n818), .A2(KEYINPUT59), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n832), .A2(KEYINPUT118), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT118), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n819), .B1(new_n830), .B2(new_n836), .ZN(G1345gat));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n277), .A3(new_n673), .ZN(new_n838));
  OAI21_X1  g637(.A(G155gat), .B1(new_n831), .B2(new_n539), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1346gat));
  INV_X1    g639(.A(new_n285), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n777), .A2(new_n841), .A3(new_n769), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT120), .Z(new_n843));
  OR2_X1    g642(.A1(new_n831), .A2(new_n599), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n285), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(G1347gat));
  NAND2_X1  g647(.A1(new_n400), .A2(new_n262), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n385), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n750), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n219), .A3(new_n609), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n468), .B1(new_n748), .B2(new_n749), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n392), .A3(new_n689), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT122), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n462), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n856), .B2(new_n219), .ZN(G1348gat));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n220), .A3(new_n572), .ZN(new_n858));
  OAI21_X1  g657(.A(G176gat), .B1(new_n851), .B2(new_n597), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1349gat));
  INV_X1    g659(.A(new_n851), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n206), .B1(new_n861), .B2(new_n673), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n854), .A2(new_n222), .A3(new_n539), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g664(.A1(new_n855), .A2(new_n207), .A3(new_n507), .ZN(new_n866));
  OAI21_X1  g665(.A(G190gat), .B1(new_n851), .B2(new_n599), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(KEYINPUT61), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(KEYINPUT61), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(G1351gat));
  NOR3_X1   g669(.A1(new_n656), .A2(new_n591), .A3(new_n359), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n853), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G197gat), .A3(new_n609), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n825), .A2(KEYINPUT123), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n821), .C1(new_n824), .C2(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n849), .A2(new_n591), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n875), .A2(new_n877), .A3(new_n462), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n879), .B2(G197gat), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT124), .ZN(G1352gat));
  NAND4_X1  g680(.A1(new_n875), .A2(new_n877), .A3(new_n572), .A4(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G204gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n872), .A2(new_n237), .A3(new_n572), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n883), .A2(new_n888), .A3(KEYINPUT126), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1353gat));
  NAND3_X1  g692(.A1(new_n872), .A2(new_n240), .A3(new_n673), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n825), .A2(new_n673), .A3(new_n878), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT63), .B1(new_n895), .B2(G211gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1354gat));
  OAI21_X1  g697(.A(new_n241), .B1(new_n873), .B2(new_n599), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n507), .A2(G218gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


