

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(KEYINPUT15), .B(n617), .Z(n943) );
  NAND2_X1 U552 ( .A1(n882), .A2(G138), .ZN(n520) );
  INV_X1 U553 ( .A(KEYINPUT95), .ZN(n657) );
  XNOR2_X1 U554 ( .A(n677), .B(n676), .ZN(n678) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n676) );
  NOR2_X1 U556 ( .A1(n675), .A2(n952), .ZN(n677) );
  NOR2_X1 U557 ( .A1(G543), .A2(n529), .ZN(n526) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NOR2_X2 U559 ( .A1(G2104), .A2(n521), .ZN(n705) );
  XNOR2_X2 U560 ( .A(n518), .B(KEYINPUT64), .ZN(n691) );
  AND2_X1 U561 ( .A1(n633), .A2(G1996), .ZN(n605) );
  XNOR2_X1 U562 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n585) );
  XNOR2_X1 U563 ( .A(n586), .B(n585), .ZN(n588) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n631) );
  XNOR2_X1 U565 ( .A(n632), .B(n631), .ZN(n639) );
  NAND2_X1 U566 ( .A1(n650), .A2(n649), .ZN(n662) );
  AND2_X1 U567 ( .A1(n731), .A2(n672), .ZN(n673) );
  NAND2_X1 U568 ( .A1(n584), .A2(n685), .ZN(n604) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n685) );
  BUF_X1 U570 ( .A(n604), .Z(n651) );
  NOR2_X1 U571 ( .A1(n733), .A2(n678), .ZN(n679) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n680) );
  INV_X1 U573 ( .A(KEYINPUT17), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n960), .A2(n682), .ZN(n725) );
  NAND2_X1 U575 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n789) );
  NOR2_X1 U577 ( .A1(G651), .A2(n565), .ZN(n790) );
  NOR2_X1 U578 ( .A1(n541), .A2(n540), .ZN(G171) );
  XNOR2_X2 U579 ( .A(n517), .B(n516), .ZN(n882) );
  INV_X1 U580 ( .A(G2105), .ZN(n521) );
  AND2_X1 U581 ( .A1(G2104), .A2(n521), .ZN(n518) );
  NAND2_X1 U582 ( .A1(G102), .A2(n691), .ZN(n519) );
  NAND2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n525) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U585 ( .A1(G114), .A2(n885), .ZN(n523) );
  NAND2_X1 U586 ( .A1(G126), .A2(n705), .ZN(n522) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(G164) );
  NAND2_X1 U589 ( .A1(G86), .A2(n789), .ZN(n528) );
  INV_X1 U590 ( .A(G651), .ZN(n529) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n526), .Z(n784) );
  NAND2_X1 U592 ( .A1(G61), .A2(n784), .ZN(n527) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n532) );
  XOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .Z(n565) );
  NOR2_X2 U595 ( .A1(n565), .A2(n529), .ZN(n785) );
  NAND2_X1 U596 ( .A1(n785), .A2(G73), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT2), .B(n530), .Z(n531) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n790), .A2(G48), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(G305) );
  NAND2_X1 U601 ( .A1(G64), .A2(n784), .ZN(n536) );
  NAND2_X1 U602 ( .A1(G52), .A2(n790), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U604 ( .A1(G77), .A2(n785), .ZN(n538) );
  NAND2_X1 U605 ( .A1(G90), .A2(n789), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NAND2_X1 U608 ( .A1(G89), .A2(n789), .ZN(n543) );
  XNOR2_X1 U609 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n785), .A2(G76), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U614 ( .A1(G63), .A2(n784), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G51), .A2(n790), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(n785), .A2(G75), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G88), .A2(n789), .ZN(n554) );
  NAND2_X1 U623 ( .A1(G62), .A2(n784), .ZN(n553) );
  NAND2_X1 U624 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U625 ( .A1(G50), .A2(n790), .ZN(n555) );
  XNOR2_X1 U626 ( .A(KEYINPUT75), .B(n555), .ZN(n556) );
  NOR2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT76), .B(n560), .Z(G166) );
  XOR2_X1 U630 ( .A(KEYINPUT82), .B(G166), .Z(G303) );
  NAND2_X1 U631 ( .A1(G49), .A2(n790), .ZN(n562) );
  NAND2_X1 U632 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U634 ( .A(KEYINPUT74), .B(n563), .ZN(n564) );
  NOR2_X1 U635 ( .A1(n784), .A2(n564), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n565), .A2(G87), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(G288) );
  NAND2_X1 U638 ( .A1(n691), .A2(G101), .ZN(n568) );
  XNOR2_X1 U639 ( .A(KEYINPUT23), .B(n568), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n882), .A2(G137), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G113), .A2(n885), .ZN(n570) );
  NAND2_X1 U642 ( .A1(G125), .A2(n705), .ZN(n569) );
  AND2_X1 U643 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n582), .A2(n580), .ZN(G160) );
  NAND2_X1 U646 ( .A1(G85), .A2(n789), .ZN(n574) );
  NAND2_X1 U647 ( .A1(G60), .A2(n784), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G72), .A2(n785), .ZN(n576) );
  NAND2_X1 U650 ( .A1(G47), .A2(n790), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(G290) );
  XNOR2_X1 U653 ( .A(G1981), .B(G305), .ZN(n960) );
  INV_X1 U654 ( .A(G40), .ZN(n579) );
  OR2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n651), .A2(G8), .ZN(n733) );
  INV_X1 U658 ( .A(n604), .ZN(n633) );
  NAND2_X1 U659 ( .A1(n633), .A2(G2072), .ZN(n586) );
  INV_X1 U660 ( .A(G1956), .ZN(n947) );
  NOR2_X1 U661 ( .A1(n633), .A2(n947), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n627) );
  NAND2_X1 U663 ( .A1(G65), .A2(n784), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G53), .A2(n790), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G78), .A2(n785), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G91), .A2(n789), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n763) );
  NAND2_X1 U670 ( .A1(n627), .A2(n763), .ZN(n626) );
  NAND2_X1 U671 ( .A1(G56), .A2(n784), .ZN(n595) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n595), .Z(n601) );
  NAND2_X1 U673 ( .A1(n789), .A2(G81), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT12), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G68), .A2(n785), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U677 ( .A(KEYINPUT13), .B(n599), .Z(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n790), .A2(G43), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n944) );
  XOR2_X1 U681 ( .A(n605), .B(KEYINPUT26), .Z(n607) );
  NAND2_X1 U682 ( .A1(n651), .A2(G1341), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n944), .A2(n608), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G92), .A2(n789), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(KEYINPUT68), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G66), .A2(n784), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G54), .A2(n790), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G79), .A2(n785), .ZN(n612) );
  XNOR2_X1 U691 ( .A(KEYINPUT69), .B(n612), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  INV_X1 U693 ( .A(n943), .ZN(n907) );
  OR2_X1 U694 ( .A1(n618), .A2(n907), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n618), .A2(n907), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G1348), .A2(n651), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n633), .A2(G2067), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n630) );
  NOR2_X1 U702 ( .A1(n627), .A2(n763), .ZN(n628) );
  XOR2_X1 U703 ( .A(n628), .B(KEYINPUT28), .Z(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n632) );
  XOR2_X1 U705 ( .A(G2078), .B(KEYINPUT25), .Z(n1005) );
  NAND2_X1 U706 ( .A1(n633), .A2(n1005), .ZN(n635) );
  NAND2_X1 U707 ( .A1(G1961), .A2(n651), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U709 ( .A(KEYINPUT90), .B(n636), .Z(n640) );
  NAND2_X1 U710 ( .A1(G171), .A2(n640), .ZN(n637) );
  XOR2_X1 U711 ( .A(KEYINPUT91), .B(n637), .Z(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n650) );
  NOR2_X1 U713 ( .A1(G171), .A2(n640), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT93), .B(n641), .Z(n646) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n733), .ZN(n664) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n651), .ZN(n661) );
  NOR2_X1 U717 ( .A1(n664), .A2(n661), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G8), .A2(n642), .ZN(n643) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n643), .ZN(n644) );
  NOR2_X1 U720 ( .A1(G168), .A2(n644), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n648) );
  XOR2_X1 U722 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n662), .A2(G286), .ZN(n656) );
  NOR2_X1 U725 ( .A1(G1971), .A2(n733), .ZN(n653) );
  NOR2_X1 U726 ( .A1(G2090), .A2(n651), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n654), .A2(G303), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n659), .A2(G8), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(KEYINPUT32), .ZN(n668) );
  NAND2_X1 U733 ( .A1(G8), .A2(n661), .ZN(n666) );
  INV_X1 U734 ( .A(n662), .ZN(n663) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n731) );
  NOR2_X1 U738 ( .A1(G1976), .A2(G288), .ZN(n949) );
  NOR2_X1 U739 ( .A1(G1971), .A2(G303), .ZN(n669) );
  XNOR2_X1 U740 ( .A(KEYINPUT96), .B(n669), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n949), .A2(n670), .ZN(n671) );
  XOR2_X1 U742 ( .A(n671), .B(KEYINPUT97), .Z(n672) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT98), .ZN(n675) );
  NAND2_X1 U744 ( .A1(G288), .A2(G1976), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(KEYINPUT99), .ZN(n952) );
  NOR2_X1 U746 ( .A1(n679), .A2(KEYINPUT33), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  INV_X1 U748 ( .A(n733), .ZN(n684) );
  AND2_X1 U749 ( .A1(KEYINPUT33), .A2(n949), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n723) );
  NAND2_X1 U751 ( .A1(G160), .A2(G40), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n687), .B(KEYINPUT83), .ZN(n750) );
  XNOR2_X1 U754 ( .A(KEYINPUT36), .B(KEYINPUT86), .ZN(n699) );
  NAND2_X1 U755 ( .A1(G116), .A2(n885), .ZN(n689) );
  NAND2_X1 U756 ( .A1(G128), .A2(n705), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n690), .B(KEYINPUT35), .ZN(n697) );
  XNOR2_X1 U759 ( .A(KEYINPUT34), .B(KEYINPUT85), .ZN(n695) );
  NAND2_X1 U760 ( .A1(G140), .A2(n882), .ZN(n693) );
  NAND2_X1 U761 ( .A1(G104), .A2(n691), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U763 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n699), .B(n698), .ZN(n901) );
  XOR2_X1 U766 ( .A(G2067), .B(KEYINPUT37), .Z(n700) );
  XNOR2_X1 U767 ( .A(KEYINPUT84), .B(n700), .ZN(n738) );
  NAND2_X1 U768 ( .A1(n901), .A2(n738), .ZN(n979) );
  NOR2_X1 U769 ( .A1(n750), .A2(n979), .ZN(n747) );
  XOR2_X1 U770 ( .A(G1986), .B(G290), .Z(n941) );
  NOR2_X1 U771 ( .A1(n941), .A2(n750), .ZN(n701) );
  NOR2_X1 U772 ( .A1(n747), .A2(n701), .ZN(n721) );
  NAND2_X1 U773 ( .A1(G131), .A2(n882), .ZN(n703) );
  NAND2_X1 U774 ( .A1(G95), .A2(n691), .ZN(n702) );
  NAND2_X1 U775 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U776 ( .A(KEYINPUT87), .B(n704), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n885), .A2(G107), .ZN(n707) );
  NAND2_X1 U778 ( .A1(G119), .A2(n705), .ZN(n706) );
  AND2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n897) );
  AND2_X1 U781 ( .A1(n897), .A2(G1991), .ZN(n719) );
  XOR2_X1 U782 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n711) );
  NAND2_X1 U783 ( .A1(G105), .A2(n691), .ZN(n710) );
  XNOR2_X1 U784 ( .A(n711), .B(n710), .ZN(n715) );
  NAND2_X1 U785 ( .A1(G129), .A2(n705), .ZN(n713) );
  NAND2_X1 U786 ( .A1(G141), .A2(n882), .ZN(n712) );
  NAND2_X1 U787 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U788 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U789 ( .A1(n885), .A2(G117), .ZN(n716) );
  NAND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n870) );
  AND2_X1 U791 ( .A1(n870), .A2(G1996), .ZN(n718) );
  NOR2_X1 U792 ( .A1(n719), .A2(n718), .ZN(n980) );
  NOR2_X1 U793 ( .A1(n980), .A2(n750), .ZN(n742) );
  INV_X1 U794 ( .A(n742), .ZN(n720) );
  NAND2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n737) );
  INV_X1 U796 ( .A(n737), .ZN(n722) );
  AND2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n755) );
  NOR2_X1 U799 ( .A1(G1981), .A2(G305), .ZN(n726) );
  XOR2_X1 U800 ( .A(n726), .B(KEYINPUT24), .Z(n727) );
  NOR2_X1 U801 ( .A1(n733), .A2(n727), .ZN(n728) );
  XNOR2_X1 U802 ( .A(KEYINPUT89), .B(n728), .ZN(n735) );
  NOR2_X1 U803 ( .A1(G2090), .A2(G303), .ZN(n729) );
  NAND2_X1 U804 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U805 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n901), .A2(n738), .ZN(n991) );
  NOR2_X1 U810 ( .A1(n870), .A2(G1996), .ZN(n739) );
  XNOR2_X1 U811 ( .A(n739), .B(KEYINPUT102), .ZN(n976) );
  NOR2_X1 U812 ( .A1(G1991), .A2(n897), .ZN(n982) );
  NOR2_X1 U813 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n982), .A2(n740), .ZN(n741) );
  NOR2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U816 ( .A1(n976), .A2(n743), .ZN(n744) );
  XNOR2_X1 U817 ( .A(n744), .B(KEYINPUT39), .ZN(n745) );
  XNOR2_X1 U818 ( .A(KEYINPUT103), .B(n745), .ZN(n746) );
  NOR2_X1 U819 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n991), .A2(n748), .ZN(n749) );
  NOR2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U822 ( .A(n751), .B(KEYINPUT104), .ZN(n752) );
  NOR2_X1 U823 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U825 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U827 ( .A(G57), .ZN(G237) );
  INV_X1 U828 ( .A(G132), .ZN(G219) );
  INV_X1 U829 ( .A(G82), .ZN(G220) );
  XOR2_X1 U830 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n758) );
  NAND2_X1 U831 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n758), .B(n757), .ZN(n759) );
  XOR2_X1 U833 ( .A(KEYINPUT65), .B(n759), .Z(n916) );
  NAND2_X1 U834 ( .A1(n916), .A2(G567), .ZN(n760) );
  XOR2_X1 U835 ( .A(KEYINPUT11), .B(n760), .Z(G234) );
  INV_X1 U836 ( .A(G860), .ZN(n766) );
  OR2_X1 U837 ( .A1(n944), .A2(n766), .ZN(G153) );
  XNOR2_X1 U838 ( .A(G171), .B(KEYINPUT67), .ZN(G301) );
  NAND2_X1 U839 ( .A1(G868), .A2(G301), .ZN(n762) );
  INV_X1 U840 ( .A(G868), .ZN(n769) );
  NAND2_X1 U841 ( .A1(n943), .A2(n769), .ZN(n761) );
  NAND2_X1 U842 ( .A1(n762), .A2(n761), .ZN(G284) );
  INV_X1 U843 ( .A(n763), .ZN(G299) );
  NOR2_X1 U844 ( .A1(G286), .A2(n769), .ZN(n765) );
  NOR2_X1 U845 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U846 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U847 ( .A1(n766), .A2(G559), .ZN(n767) );
  NAND2_X1 U848 ( .A1(n767), .A2(n907), .ZN(n768) );
  XNOR2_X1 U849 ( .A(n768), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U850 ( .A1(G559), .A2(n769), .ZN(n770) );
  NAND2_X1 U851 ( .A1(n907), .A2(n770), .ZN(n771) );
  XNOR2_X1 U852 ( .A(n771), .B(KEYINPUT71), .ZN(n773) );
  NOR2_X1 U853 ( .A1(n944), .A2(G868), .ZN(n772) );
  NOR2_X1 U854 ( .A1(n773), .A2(n772), .ZN(G282) );
  NAND2_X1 U855 ( .A1(n705), .A2(G123), .ZN(n774) );
  XNOR2_X1 U856 ( .A(n774), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U857 ( .A1(G135), .A2(n882), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U859 ( .A(KEYINPUT72), .B(n777), .ZN(n781) );
  NAND2_X1 U860 ( .A1(G111), .A2(n885), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G99), .A2(n691), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U863 ( .A1(n781), .A2(n780), .ZN(n981) );
  XNOR2_X1 U864 ( .A(G2096), .B(n981), .ZN(n782) );
  INV_X1 U865 ( .A(G2100), .ZN(n847) );
  NAND2_X1 U866 ( .A1(n782), .A2(n847), .ZN(G156) );
  NAND2_X1 U867 ( .A1(n907), .A2(G559), .ZN(n806) );
  XNOR2_X1 U868 ( .A(n944), .B(n806), .ZN(n783) );
  NOR2_X1 U869 ( .A1(n783), .A2(G860), .ZN(n795) );
  NAND2_X1 U870 ( .A1(n784), .A2(G67), .ZN(n788) );
  NAND2_X1 U871 ( .A1(G80), .A2(n785), .ZN(n786) );
  XOR2_X1 U872 ( .A(KEYINPUT73), .B(n786), .Z(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n794) );
  NAND2_X1 U874 ( .A1(G93), .A2(n789), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G55), .A2(n790), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n797) );
  XNOR2_X1 U878 ( .A(n795), .B(n797), .ZN(G145) );
  NOR2_X1 U879 ( .A1(G868), .A2(n797), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(KEYINPUT79), .ZN(n809) );
  XNOR2_X1 U881 ( .A(G305), .B(G290), .ZN(n805) );
  XNOR2_X1 U882 ( .A(n944), .B(G288), .ZN(n803) );
  XNOR2_X1 U883 ( .A(KEYINPUT19), .B(KEYINPUT77), .ZN(n799) );
  XOR2_X1 U884 ( .A(n797), .B(KEYINPUT78), .Z(n798) );
  XNOR2_X1 U885 ( .A(n799), .B(n798), .ZN(n800) );
  XOR2_X1 U886 ( .A(G299), .B(n800), .Z(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(G166), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n805), .B(n804), .ZN(n904) );
  XNOR2_X1 U890 ( .A(n904), .B(n806), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G868), .A2(n807), .ZN(n808) );
  NAND2_X1 U892 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2084), .A2(G2078), .ZN(n810) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U895 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U898 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U899 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U901 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U902 ( .A1(G96), .A2(n816), .ZN(n839) );
  NAND2_X1 U903 ( .A1(G2106), .A2(n839), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n817), .B(KEYINPUT80), .ZN(n821) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U906 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U907 ( .A1(G108), .A2(n819), .ZN(n840) );
  NAND2_X1 U908 ( .A1(G567), .A2(n840), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U910 ( .A(KEYINPUT81), .B(n822), .Z(n841) );
  NAND2_X1 U911 ( .A1(G661), .A2(G483), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n841), .A2(n823), .ZN(n838) );
  NAND2_X1 U913 ( .A1(n838), .A2(G36), .ZN(G176) );
  XNOR2_X1 U914 ( .A(G2435), .B(G2451), .ZN(n833) );
  XOR2_X1 U915 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n825) );
  XNOR2_X1 U916 ( .A(G2454), .B(G2430), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U918 ( .A(G2446), .B(G2438), .Z(n827) );
  XNOR2_X1 U919 ( .A(G1348), .B(G1341), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U921 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U922 ( .A(G2427), .B(G2443), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U925 ( .A1(n834), .A2(G14), .ZN(n910) );
  XNOR2_X1 U926 ( .A(KEYINPUT107), .B(n910), .ZN(G401) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n916), .ZN(G217) );
  NAND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  XOR2_X1 U929 ( .A(KEYINPUT108), .B(n835), .Z(n836) );
  NAND2_X1 U930 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n841), .ZN(G319) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2067), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(G2096), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n851) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2678), .Z(n849) );
  XOR2_X1 U947 ( .A(KEYINPUT109), .B(n847), .Z(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(G227) );
  XOR2_X1 U950 ( .A(KEYINPUT110), .B(G1991), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1996), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U953 ( .A(n854), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1971), .B(G1976), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(G1986), .B(G1981), .Z(n858) );
  XOR2_X1 U957 ( .A(G1966), .B(n947), .Z(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U960 ( .A(KEYINPUT111), .B(G2474), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G124), .A2(n705), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n885), .A2(G112), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G136), .A2(n882), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G100), .A2(n691), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U970 ( .A(G160), .B(n870), .Z(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(n981), .ZN(n881) );
  NAND2_X1 U972 ( .A1(G142), .A2(n882), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G106), .A2(n691), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT45), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G118), .A2(n885), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n705), .A2(G130), .ZN(n877) );
  XOR2_X1 U979 ( .A(KEYINPUT112), .B(n877), .Z(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(n881), .B(n880), .Z(n892) );
  NAND2_X1 U982 ( .A1(G139), .A2(n882), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G103), .A2(n691), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n890) );
  NAND2_X1 U985 ( .A1(G115), .A2(n885), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G127), .A2(n705), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n969) );
  XNOR2_X1 U990 ( .A(n969), .B(G162), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n894) );
  XNOR2_X1 U993 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(n896), .B(n895), .Z(n899) );
  XOR2_X1 U996 ( .A(G164), .B(n897), .Z(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(n903) );
  XOR2_X1 U1000 ( .A(KEYINPUT115), .B(n903), .Z(G395) );
  XNOR2_X1 U1001 ( .A(n904), .B(KEYINPUT116), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(G171), .B(G286), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n909), .ZN(G397) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n910), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n916), .ZN(G223) );
  XNOR2_X1 U1015 ( .A(G1348), .B(KEYINPUT59), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n917), .B(G4), .ZN(n921) );
  XOR2_X1 U1017 ( .A(n947), .B(G20), .Z(n919) );
  XNOR2_X1 U1018 ( .A(G6), .B(G1981), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1021 ( .A(KEYINPUT127), .B(G1341), .Z(n922) );
  XNOR2_X1 U1022 ( .A(G19), .B(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT60), .B(n925), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G21), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(G5), .B(G1961), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G22), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(G24), .B(G1986), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G1976), .B(G23), .Z(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT61), .B(n937), .ZN(n938) );
  INV_X1 U1037 ( .A(G16), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n940), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n939), .A2(G11), .ZN(n968) );
  XOR2_X1 U1040 ( .A(KEYINPUT56), .B(n940), .Z(n965) );
  XNOR2_X1 U1041 ( .A(G171), .B(G1961), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n958) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n943), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(n944), .B(G1341), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G299), .B(n947), .Z(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1048 ( .A(G1971), .B(G303), .Z(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1051 ( .A(KEYINPUT125), .B(n954), .Z(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G168), .B(G1966), .Z(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1056 ( .A(KEYINPUT57), .B(n961), .Z(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1059 ( .A(KEYINPUT126), .B(n966), .Z(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n1001) );
  XOR2_X1 U1061 ( .A(G2072), .B(n969), .Z(n971) );
  XOR2_X1 U1062 ( .A(G164), .B(G2078), .Z(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT50), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n974), .B(n973), .ZN(n994) );
  XOR2_X1 U1067 ( .A(G2090), .B(G162), .Z(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT51), .B(n977), .Z(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT118), .B(n978), .ZN(n989) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n987) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1073 ( .A(G160), .B(G2084), .Z(n983) );
  XNOR2_X1 U1074 ( .A(KEYINPUT117), .B(n983), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(KEYINPUT119), .B(n992), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1081 ( .A(n995), .B(KEYINPUT52), .Z(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n996), .ZN(n997) );
  NOR2_X1 U1083 ( .A1(KEYINPUT55), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT123), .B(n998), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n999), .A2(G29), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1022) );
  XOR2_X1 U1087 ( .A(G2090), .B(G35), .Z(n1015) );
  XOR2_X1 U1088 ( .A(G25), .B(G1991), .Z(n1002) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(G28), .ZN(n1011) );
  XNOR2_X1 U1090 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G33), .B(G2072), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(n1005), .B(G27), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1996), .B(G32), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(KEYINPUT53), .B(n1012), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT124), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(KEYINPUT54), .B(G2084), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G34), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT55), .B(n1019), .Z(n1020) );
  NOR2_X1 U1105 ( .A1(G29), .A2(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(n1023), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

