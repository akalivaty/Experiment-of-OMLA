//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT66), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G2104), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(new_n466), .A3(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n459), .A2(new_n460), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT64), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G125), .C1(new_n471), .C2(new_n472), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(G2105), .B2(new_n478), .ZN(G160));
  AND2_X1   g054(.A1(new_n461), .A2(new_n466), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n461), .A2(new_n466), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT68), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n484), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT69), .Z(new_n491));
  NAND2_X1  g066(.A1(new_n480), .A2(new_n484), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(G136), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n461), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(G2104), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n497), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n498), .B1(new_n497), .B2(new_n505), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT4), .A2(G138), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n461), .A2(new_n466), .A3(new_n484), .A4(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(G138), .B(new_n484), .C1(new_n471), .C2(new_n472), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(G164));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  INV_X1    g096(.A(new_n517), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n523), .B1(new_n518), .B2(KEYINPUT72), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n520), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  INV_X1    g112(.A(new_n527), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n517), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n536), .A2(new_n537), .B1(G89), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n519), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT74), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n519), .A2(G52), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G90), .Z(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n531), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT76), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(KEYINPUT76), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G651), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n539), .A2(G81), .B1(G43), .B2(new_n519), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT78), .Z(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT79), .Z(G188));
  AOI22_X1  g143(.A1(new_n527), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n531), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n539), .A2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n519), .A2(G53), .ZN(new_n572));
  NOR2_X1   g147(.A1(KEYINPUT80), .A2(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g149(.A(KEYINPUT80), .B(KEYINPUT9), .Z(new_n575));
  NAND3_X1  g150(.A1(new_n519), .A2(G53), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n570), .A2(new_n571), .A3(new_n574), .A4(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n539), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n519), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n538), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n519), .A2(G48), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n528), .A2(KEYINPUT81), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT81), .B1(new_n528), .B2(new_n590), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n539), .A2(G85), .B1(G47), .B2(new_n519), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n531), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n519), .A2(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n519), .A2(KEYINPUT82), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n600), .A2(G54), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OR3_X1    g178(.A1(new_n528), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n527), .A2(G66), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT83), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT10), .B1(new_n528), .B2(new_n603), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n602), .A2(new_n604), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n599), .B1(new_n611), .B2(G868), .ZN(G321));
  XOR2_X1   g187(.A(G321), .B(KEYINPUT84), .Z(G284));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G299), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT85), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n559), .ZN(G323));
  XOR2_X1   g198(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  AOI22_X1  g200(.A1(new_n486), .A2(G123), .B1(G135), .B2(new_n493), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n484), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  OR2_X1    g205(.A1(new_n471), .A2(new_n472), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(new_n484), .A3(new_n468), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT88), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n648), .B2(new_n649), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT88), .B1(new_n648), .B2(new_n649), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT89), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT90), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n660), .B(KEYINPUT17), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n658), .A3(new_n661), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT92), .Z(new_n667));
  INV_X1    g242(.A(new_n661), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n659), .B2(new_n660), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT91), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n658), .B2(new_n665), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2096), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n636), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT93), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n682), .A2(new_n683), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n679), .A2(new_n684), .A3(new_n681), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(new_n683), .C2(new_n682), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT22), .B(G1981), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G2090), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n495), .A2(G29), .ZN(new_n696));
  INV_X1    g271(.A(G35), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(G29), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n696), .B(new_n700), .C1(G29), .C2(new_n697), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n695), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT31), .B(G11), .Z(new_n703));
  OR2_X1    g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(KEYINPUT24), .A2(G34), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G160), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2084), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  NAND2_X1  g285(.A1(G171), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G5), .B2(G16), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n703), .B(new_n709), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(G29), .A2(G33), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n631), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(new_n484), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT100), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n493), .A2(G139), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(new_n705), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2072), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n626), .A2(G29), .A3(new_n628), .ZN(new_n724));
  NAND2_X1  g299(.A1(G299), .A2(G16), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n726), .A2(KEYINPUT23), .A3(G20), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT23), .ZN(new_n728));
  INV_X1    g303(.A(G20), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G16), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n725), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1956), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT30), .B(G28), .Z(new_n733));
  OAI22_X1  g308(.A1(new_n712), .A2(new_n710), .B1(G29), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n713), .A2(new_n723), .A3(new_n724), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n726), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n726), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1966), .ZN(new_n739));
  OR3_X1    g314(.A1(new_n702), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(G4), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n611), .B2(new_n726), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT97), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT96), .B(G1348), .Z(new_n744));
  XOR2_X1   g319(.A(new_n743), .B(new_n744), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n726), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n559), .B2(new_n726), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1341), .Z(new_n748));
  INV_X1    g323(.A(G26), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(G29), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT28), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n486), .A2(G128), .B1(G140), .B2(new_n493), .ZN(new_n753));
  NOR2_X1   g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(new_n484), .B2(G116), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n752), .B1(new_n756), .B2(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n751), .A2(KEYINPUT28), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT98), .B(G2067), .Z(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n745), .A2(new_n748), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n745), .A2(KEYINPUT99), .A3(new_n748), .A4(new_n762), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n740), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G23), .ZN(new_n768));
  AND3_X1   g343(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(G288), .A2(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n726), .A2(G6), .ZN(new_n777));
  INV_X1    g352(.A(G305), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n726), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1981), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n726), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n726), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n776), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n776), .A2(new_n782), .A3(KEYINPUT34), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n486), .A2(G119), .B1(G131), .B2(new_n493), .ZN(new_n792));
  NOR2_X1   g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(new_n484), .B2(G107), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  MUX2_X1   g374(.A(G24), .B(G290), .S(G16), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1986), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n791), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT36), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n791), .A2(new_n805), .A3(new_n802), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n699), .A2(new_n695), .A3(new_n701), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT102), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n705), .A2(G27), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G164), .B2(new_n705), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n767), .A2(new_n807), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n486), .A2(G129), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G2105), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT101), .B(KEYINPUT26), .Z(new_n818));
  NAND3_X1  g393(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G29), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G29), .B2(G32), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT27), .B(G1996), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n814), .A2(new_n826), .ZN(G311));
  AND3_X1   g402(.A1(new_n767), .A2(new_n807), .A3(new_n809), .ZN(new_n828));
  INV_X1    g403(.A(new_n826), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n828), .A2(KEYINPUT103), .A3(new_n829), .A4(new_n813), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n814), .B2(new_n826), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G150));
  AOI22_X1  g408(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT104), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G651), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n539), .A2(G93), .B1(G55), .B2(new_n519), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n559), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n558), .A2(new_n837), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n611), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT105), .ZN(new_n846));
  AOI21_X1  g421(.A(G860), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n838), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(G145));
  XOR2_X1   g426(.A(new_n721), .B(new_n756), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n486), .A2(G130), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n493), .A2(G142), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n484), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT106), .Z(new_n857));
  OAI211_X1 g432(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n509), .A2(new_n497), .A3(new_n512), .A4(new_n505), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n634), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n795), .B(new_n821), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n629), .B(G160), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n495), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n495), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n865), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n873), .A2(new_n862), .A3(new_n869), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n860), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n862), .B1(new_n873), .B2(new_n869), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n863), .A3(new_n871), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n859), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g456(.A(new_n621), .B(new_n841), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n610), .A2(G299), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n610), .A2(G299), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(KEYINPUT41), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n887), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n773), .A2(KEYINPUT107), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n773), .A2(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G166), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n778), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n778), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n902), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n906), .A2(new_n898), .A3(new_n899), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n905), .A2(new_n907), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n894), .A2(new_n910), .A3(new_n896), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n911), .A3(G868), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT108), .B1(new_n838), .B2(new_n614), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT108), .A4(G868), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(G295));
  AND2_X1   g491(.A1(new_n914), .A2(new_n915), .ZN(G331));
  INV_X1    g492(.A(new_n886), .ZN(new_n918));
  NAND2_X1  g493(.A1(G168), .A2(G301), .ZN(new_n919));
  NAND2_X1  g494(.A1(G286), .A2(G171), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n841), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n919), .A2(new_n839), .A3(new_n840), .A4(new_n920), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT109), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(KEYINPUT109), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n891), .B1(new_n922), .B2(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n908), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n890), .A4(new_n888), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n922), .A2(new_n886), .A3(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n910), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n931), .A3(new_n876), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n932), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n930), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n908), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n876), .A3(new_n931), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n939), .B2(KEYINPUT43), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n935), .A2(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n932), .A2(KEYINPUT112), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n928), .A2(new_n931), .A3(new_n948), .A4(new_n876), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(KEYINPUT43), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n950), .A3(KEYINPUT44), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(G397));
  NAND2_X1  g530(.A1(new_n467), .A2(new_n469), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n484), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n478), .A2(G2105), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(G40), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT45), .B1(new_n861), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n756), .B(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(new_n822), .ZN(new_n968));
  OAI221_X1 g543(.A(new_n965), .B1(KEYINPUT126), .B2(KEYINPUT46), .C1(new_n968), .C2(new_n962), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n822), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n821), .A2(G1996), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n795), .A2(new_n797), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n974), .A2(new_n976), .B1(G2067), .B2(new_n756), .ZN(new_n977));
  INV_X1    g552(.A(new_n962), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n795), .A2(new_n797), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n974), .A2(new_n984), .A3(new_n975), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n985), .B2(new_n962), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n970), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT115), .B(G1981), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n589), .A2(new_n593), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n587), .A2(new_n588), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n528), .A2(new_n590), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n957), .A2(new_n958), .A3(G40), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n861), .A2(new_n960), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n989), .A2(new_n992), .A3(KEYINPUT49), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n771), .B2(new_n772), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1003), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1000), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1000), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1002), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n509), .A2(new_n512), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n497), .A2(new_n505), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n996), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(new_n695), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n497), .A2(new_n505), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT71), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n497), .A2(new_n498), .A3(new_n505), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n1021), .B2(new_n960), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n1023));
  NAND3_X1  g598(.A1(G160), .A2(new_n1023), .A3(G40), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n785), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n999), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G166), .A2(new_n999), .ZN(new_n1027));
  AND2_X1   g602(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1028));
  NOR2_X1   g603(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1010), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n959), .B(new_n1034), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1021), .A2(new_n1015), .A3(new_n960), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n957), .A2(new_n958), .A3(new_n1015), .A4(G40), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(KEYINPUT116), .C1(new_n996), .C2(new_n997), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1025), .B1(new_n1039), .B2(G2090), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1031), .B1(new_n1040), .B2(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT123), .B(G1961), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1015), .B1(new_n1021), .B2(new_n960), .ZN(new_n1044));
  OAI211_X1 g619(.A(G160), .B(G40), .C1(new_n997), .C2(KEYINPUT50), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n961), .A2(new_n996), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2078), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1021), .A2(new_n960), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1047), .B(new_n1049), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1022), .A2(new_n1024), .A3(G2078), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1046), .B(new_n1052), .C1(new_n1053), .C2(KEYINPUT53), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G301), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(new_n1023), .A3(new_n1049), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1046), .B(new_n1056), .C1(new_n1053), .C2(KEYINPUT53), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1055), .B(KEYINPUT54), .C1(G301), .C2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT124), .B1(new_n1057), .B2(G171), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(G171), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n996), .B1(new_n1014), .B2(KEYINPUT45), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n812), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1048), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(G301), .A3(new_n1046), .A4(new_n1056), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(KEYINPUT124), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1058), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G2084), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1011), .A2(new_n1070), .A3(new_n1016), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1011), .A2(new_n1016), .A3(KEYINPUT117), .A4(new_n1070), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1073), .A2(G168), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(G286), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1069), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(G299), .B(KEYINPUT57), .ZN(new_n1086));
  INV_X1    g661(.A(G1956), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1039), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT120), .B(G2072), .Z(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT56), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1063), .A2(new_n1064), .A3(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1088), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1089), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1086), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1086), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1088), .A2(new_n1096), .A3(new_n1092), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1063), .A2(new_n971), .A3(new_n1064), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n996), .B2(new_n997), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n558), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1088), .A2(new_n1096), .A3(new_n1092), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1096), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1014), .A2(G160), .A3(G40), .A4(new_n966), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n998), .A2(KEYINPUT121), .A3(new_n966), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1348), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n610), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1115), .A4(new_n611), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1098), .A2(new_n1104), .A3(new_n1108), .A4(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n610), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1095), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1085), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1083), .A2(new_n1079), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1081), .B1(new_n1078), .B2(G8), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT62), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1060), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1080), .B(new_n1131), .C1(new_n1079), .C2(new_n1083), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1042), .B1(new_n1126), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1010), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n1032), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1002), .A2(new_n1003), .A3(new_n769), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n989), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1000), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT63), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1082), .A2(new_n1142), .A3(G8), .A4(G168), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1082), .A2(G8), .A3(G168), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT118), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1141), .B(new_n1033), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1143), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1042), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1140), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1135), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n985), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(G1986), .B2(G290), .ZN(new_n1154));
  INV_X1    g729(.A(new_n980), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n962), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT125), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1108), .A2(new_n1120), .A3(new_n1104), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1124), .B1(new_n1159), .B2(new_n1098), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1133), .B1(new_n1160), .B2(new_n1085), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1150), .B1(new_n1161), .B2(new_n1042), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1162), .A2(new_n1163), .A3(new_n1156), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n987), .B1(new_n1158), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g740(.A1(new_n880), .A2(new_n656), .A3(new_n674), .ZN(new_n1167));
  NAND4_X1  g741(.A1(new_n1167), .A2(new_n943), .A3(G319), .A4(new_n693), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


