//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n448, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(new_n442), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n460), .A2(new_n457), .B1(new_n455), .B2(new_n451), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n469), .A2(KEYINPUT70), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT70), .B1(new_n469), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n464), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT71), .B(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n478), .A2(new_n480), .B1(new_n481), .B2(G101), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n475), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n478), .A2(new_n472), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT73), .Z(new_n489));
  OR2_X1    g064(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI221_X1 g067(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n492), .C2(G112), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT74), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT3), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n464), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(G136), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  INV_X1    g077(.A(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(G102), .A3(G2104), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT3), .B(G2104), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n492), .A2(new_n506), .A3(G138), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n490), .B2(new_n491), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n511), .A2(new_n497), .A3(KEYINPUT4), .A4(new_n464), .ZN(new_n512));
  NAND2_X1  g087(.A1(G114), .A2(G2104), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n478), .B2(G126), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n509), .B(new_n512), .C1(new_n515), .C2(new_n503), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT77), .B1(new_n518), .B2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(G543), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(new_n522), .B1(KEYINPUT5), .B2(new_n518), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(KEYINPUT6), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(KEYINPUT76), .A3(G651), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT75), .B1(new_n527), .B2(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(new_n525), .A3(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n523), .A2(new_n529), .A3(G88), .A4(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G50), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n533), .A2(G543), .A3(new_n526), .A4(new_n528), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(G75), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n523), .B2(G62), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n525), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G166));
  NAND2_X1  g116(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n529), .A2(new_n543), .A3(G543), .A4(new_n533), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n529), .A2(G89), .A3(new_n533), .ZN(new_n547));
  NAND2_X1  g122(.A1(G63), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(new_n523), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n551));
  NAND3_X1  g126(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n546), .A2(new_n550), .A3(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n542), .B2(new_n544), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n525), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n523), .A2(new_n529), .A3(new_n533), .ZN(new_n562));
  INV_X1    g137(.A(G90), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n558), .A2(new_n561), .A3(new_n565), .ZN(G301));
  INV_X1    g141(.A(G301), .ZN(G171));
  INV_X1    g142(.A(G43), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n542), .B2(new_n544), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n525), .ZN(new_n571));
  INV_X1    g146(.A(G81), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  NOR3_X1   g148(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  AND3_X1   g150(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G36), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G188));
  AOI22_X1  g155(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n525), .ZN(new_n582));
  INV_X1    g157(.A(new_n562), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n582), .B1(G91), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(G53), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n536), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n536), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(KEYINPUT9), .A3(G53), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n584), .A2(new_n587), .A3(new_n589), .ZN(G299));
  AND2_X1   g165(.A1(new_n523), .A2(G62), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n591), .B2(new_n538), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(G50), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n592), .A2(KEYINPUT80), .A3(new_n534), .A4(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n537), .B2(new_n540), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G303));
  NAND2_X1  g172(.A1(new_n583), .A2(G87), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n588), .A2(G49), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G288));
  AOI22_X1  g176(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n525), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n583), .A2(G86), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n588), .A2(G48), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n545), .A2(G47), .B1(new_n583), .B2(G85), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT81), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n525), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n523), .A2(new_n529), .A3(G92), .A4(new_n533), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT10), .Z(new_n613));
  AOI22_X1  g188(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n525), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G54), .B2(new_n545), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n613), .A2(new_n616), .A3(KEYINPUT82), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT82), .B1(new_n613), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(new_n619), .B2(G868), .ZN(G284));
  XOR2_X1   g195(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n589), .A2(new_n587), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n583), .A2(G91), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n623), .A2(new_n624), .A3(new_n582), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n622), .B1(G868), .B2(new_n625), .ZN(G297));
  OAI21_X1  g201(.A(new_n622), .B1(G868), .B2(new_n625), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n619), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n619), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n574), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g208(.A1(new_n487), .A2(G123), .B1(G135), .B2(new_n499), .ZN(new_n634));
  OAI221_X1 g209(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n492), .C2(G111), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n481), .A2(new_n506), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2451), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT85), .Z(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT17), .Z(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n659), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n669), .B2(new_n659), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2096), .Z(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2100), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n687), .C1(new_n685), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(G1986), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G1981), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n487), .A2(G119), .B1(G131), .B2(new_n499), .ZN(new_n698));
  OAI221_X1 g273(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n492), .C2(G107), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n697), .B1(new_n700), .B2(new_n696), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G24), .B(G290), .S(G16), .Z(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G6), .B(G305), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT87), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G23), .ZN(new_n716));
  INV_X1    g291(.A(G288), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT33), .B(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n710), .A2(new_n715), .A3(new_n720), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n703), .B(new_n706), .C1(new_n721), .C2(KEYINPUT34), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT88), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n723), .A2(new_n727), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n696), .A2(G35), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n501), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g308(.A1(G160), .A2(G29), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G34), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(new_n737), .A3(new_n696), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT26), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n487), .B2(G129), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G105), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n499), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G29), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n741), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(G171), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G5), .B2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n730), .A2(new_n733), .B1(new_n756), .B2(KEYINPUT92), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n711), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n619), .B2(new_n711), .ZN(new_n759));
  INV_X1    g334(.A(G1348), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n733), .A2(new_n730), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n711), .A2(KEYINPUT23), .A3(G20), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n764));
  INV_X1    g339(.A(G20), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G16), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n766), .C1(new_n625), .C2(new_n711), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT93), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n729), .A2(new_n757), .A3(new_n761), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G168), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G16), .B2(G21), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n696), .A2(G26), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n487), .A2(G128), .B1(G140), .B2(new_n499), .ZN(new_n776));
  OAI221_X1 g351(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n492), .C2(G116), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n775), .B1(new_n779), .B2(new_n696), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n775), .B(new_n780), .S(KEYINPUT28), .Z(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n762), .A2(KEYINPUT93), .A3(new_n768), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n711), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n574), .B2(new_n711), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT89), .B(G1341), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G29), .B2(G33), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n791), .A2(G29), .A3(G33), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n492), .A2(G103), .A3(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT91), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT25), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n506), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n492), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G139), .B2(new_n499), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n792), .B(new_n793), .C1(new_n802), .C2(new_n696), .ZN(new_n803));
  INV_X1    g378(.A(G2072), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n772), .A2(new_n773), .ZN(new_n806));
  NOR2_X1   g381(.A1(G27), .A2(G29), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G164), .B2(G29), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G2078), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n739), .A2(new_n740), .ZN(new_n812));
  AOI211_X1 g387(.A(new_n811), .B(new_n812), .C1(new_n803), .C2(new_n804), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT30), .B(G28), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n750), .A2(new_n751), .B1(new_n696), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n813), .B(new_n815), .C1(G2078), .C2(new_n808), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n756), .A2(KEYINPUT92), .B1(new_n753), .B2(new_n755), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n636), .A2(new_n696), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n790), .A2(new_n805), .A3(new_n806), .A4(new_n819), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n770), .A2(new_n774), .A3(new_n784), .A4(new_n820), .ZN(G311));
  NOR2_X1   g396(.A1(new_n770), .A2(new_n820), .ZN(new_n822));
  INV_X1    g397(.A(new_n774), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(new_n823), .A3(new_n783), .ZN(G150));
  XOR2_X1   g399(.A(KEYINPUT94), .B(G55), .Z(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n542), .B2(new_n544), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n827), .A2(new_n525), .B1(new_n562), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n574), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n545), .A2(G43), .ZN(new_n833));
  INV_X1    g408(.A(new_n571), .ZN(new_n834));
  INV_X1    g409(.A(new_n573), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n830), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n619), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT95), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n830), .A2(new_n843), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n778), .B(G164), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(new_n748), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n748), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n801), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n802), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n499), .A2(G142), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT97), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n487), .A2(G130), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT98), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(G118), .B2(new_n492), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n639), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n700), .Z(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n501), .B(new_n636), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G160), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n856), .A2(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n856), .A2(new_n865), .ZN(new_n873));
  INV_X1    g448(.A(new_n865), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n854), .A2(new_n874), .A3(new_n855), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n869), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g453(.A(KEYINPUT99), .B(new_n869), .C1(new_n873), .C2(new_n875), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n871), .B(new_n872), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g456(.A1(G299), .A2(new_n616), .A3(new_n613), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n613), .A2(new_n616), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n625), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT101), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(KEYINPUT101), .B2(new_n882), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n887), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n832), .A2(new_n837), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n630), .B(new_n892), .ZN(new_n893));
  MUX2_X1   g468(.A(new_n891), .B(new_n890), .S(new_n893), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT42), .ZN(new_n895));
  XOR2_X1   g470(.A(G288), .B(G166), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G305), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(G290), .Z(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT102), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n895), .B(new_n900), .ZN(new_n901));
  MUX2_X1   g476(.A(new_n831), .B(new_n901), .S(G868), .Z(G295));
  MUX2_X1   g477(.A(new_n831), .B(new_n901), .S(G868), .Z(G331));
  NAND2_X1  g478(.A1(new_n885), .A2(KEYINPUT41), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n889), .A2(new_n886), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n557), .A2(new_n564), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n561), .ZN(new_n908));
  NOR4_X1   g483(.A1(new_n557), .A2(new_n560), .A3(new_n564), .A4(KEYINPUT103), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(G286), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(G301), .A2(KEYINPUT103), .A3(G286), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n892), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G301), .A2(KEYINPUT103), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n906), .A3(new_n561), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(G168), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n838), .A3(new_n911), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT104), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(KEYINPUT104), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n904), .B(new_n905), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT105), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n916), .A2(new_n838), .A3(new_n911), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n838), .B1(new_n916), .B2(new_n911), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n919), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n904), .A4(new_n905), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n890), .A2(new_n917), .A3(new_n913), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n922), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n931), .A2(KEYINPUT106), .A3(new_n898), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n931), .B2(new_n898), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n891), .B1(new_n924), .B2(new_n925), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n890), .A3(new_n919), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n872), .B1(new_n937), .B2(new_n898), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n938), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(new_n937), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n940), .B(new_n941), .C1(new_n899), .C2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n941), .B(new_n940), .C1(new_n932), .C2(new_n933), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n942), .A2(new_n899), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n947), .B2(new_n938), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI211_X1 g526(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n946), .C2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  OAI21_X1  g529(.A(G138), .B1(new_n470), .B2(new_n471), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n464), .A2(new_n466), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n508), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n512), .A2(new_n957), .A3(new_n504), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n497), .A2(G126), .A3(new_n464), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n503), .B1(new_n959), .B2(new_n513), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n954), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT108), .B(G40), .Z(new_n964));
  OAI211_X1 g539(.A(new_n482), .B(new_n964), .C1(new_n473), .C2(new_n474), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n778), .B(G2067), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(new_n747), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n963), .A2(G1996), .A3(new_n965), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n969), .B(new_n971), .Z(new_n972));
  OAI211_X1 g547(.A(new_n968), .B(new_n972), .C1(KEYINPUT126), .C2(new_n970), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT47), .Z(new_n974));
  NOR2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n966), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT48), .Z(new_n977));
  XNOR2_X1  g552(.A(new_n700), .B(new_n702), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT109), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n747), .B(G1996), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(new_n967), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n982), .B2(new_n966), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n700), .A2(new_n702), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT125), .Z(new_n985));
  OAI22_X1  g560(.A1(new_n985), .A2(new_n981), .B1(G2067), .B2(new_n778), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n974), .B(new_n983), .C1(new_n966), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n965), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n954), .C1(new_n958), .C2(new_n960), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n963), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n714), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT50), .B1(new_n516), .B2(new_n954), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT50), .B(new_n954), .C1(new_n958), .C2(new_n960), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n730), .B(new_n988), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n991), .B2(new_n995), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(G303), .B2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  AOI211_X1 g577(.A(KEYINPUT55), .B(new_n1002), .C1(new_n594), .C2(new_n596), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n999), .A2(KEYINPUT111), .A3(G8), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n991), .A2(new_n995), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(G8), .A3(new_n1004), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1004), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n965), .A2(new_n961), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(new_n1002), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n717), .A2(G1976), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(KEYINPUT52), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT113), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(G305), .A2(G1981), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(G305), .B2(G1981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1028), .A2(new_n1031), .A3(new_n1029), .A4(KEYINPUT49), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1025), .A2(new_n1027), .B1(new_n1036), .B2(new_n1017), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n961), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n965), .B1(new_n1039), .B2(new_n993), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n740), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n990), .A2(new_n773), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(G168), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G286), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1012), .A2(new_n1015), .A3(new_n1037), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT63), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(KEYINPUT116), .A3(new_n1047), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n999), .A2(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1047), .B1(new_n1052), .B2(new_n1013), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1012), .A2(new_n1053), .A3(new_n1037), .A4(new_n1045), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT117), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1012), .A2(new_n1037), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1045), .A4(new_n1053), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1050), .A2(new_n1051), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1037), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1034), .A2(new_n1017), .A3(new_n1035), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1022), .A3(new_n717), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1028), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1017), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT115), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1059), .A2(new_n1060), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1060), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1056), .A2(new_n1015), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G299), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n625), .A2(KEYINPUT57), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n990), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1074), .B(new_n1077), .C1(G1956), .C2(new_n1040), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1040), .A2(KEYINPUT119), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1040), .A2(KEYINPUT119), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(G1348), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1016), .A2(new_n782), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1078), .B(new_n619), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1040), .A2(G1956), .B1(new_n990), .B2(new_n1076), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n990), .A2(KEYINPUT121), .A3(G1996), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT121), .B1(new_n990), .B2(G1996), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT58), .B(G1341), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1016), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n574), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT59), .ZN(new_n1096));
  INV_X1    g671(.A(new_n619), .ZN(new_n1097));
  OR4_X1    g672(.A1(KEYINPUT60), .A2(new_n1081), .A3(new_n1097), .A4(new_n1083), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1040), .B(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n760), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1101), .B2(new_n1082), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1081), .A2(new_n619), .A3(new_n1083), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1078), .A2(new_n1086), .A3(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT61), .B1(new_n1078), .B2(new_n1086), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1096), .A2(new_n1098), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1089), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1100), .A2(new_n753), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n990), .A2(G2078), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1119), .A3(G171), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1100), .A2(new_n753), .B1(new_n1113), .B2(new_n1112), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  OAI21_X1  g698(.A(G40), .B1(new_n483), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(G2078), .B(new_n1124), .C1(new_n1123), .C2(new_n483), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1113), .B1(new_n469), .B2(new_n472), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n963), .A3(new_n989), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1110), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(G171), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1111), .A2(G301), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(KEYINPUT54), .ZN(new_n1135));
  AOI21_X1  g710(.A(G301), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1044), .A2(KEYINPUT51), .ZN(new_n1139));
  AOI21_X1  g714(.A(G168), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT51), .ZN(new_n1141));
  OAI211_X1 g716(.A(G8), .B(new_n1043), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1109), .A2(new_n1130), .A3(new_n1138), .A4(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1139), .A2(new_n1142), .A3(KEYINPUT62), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT62), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1121), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1070), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1068), .A2(new_n1069), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n982), .ZN(new_n1150));
  XNOR2_X1  g725(.A(G290), .B(new_n705), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n963), .B(new_n965), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n987), .B1(new_n1149), .B2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g728(.A1(new_n674), .A2(new_n656), .A3(G319), .ZN(new_n1155));
  XOR2_X1   g729(.A(new_n1155), .B(KEYINPUT127), .Z(new_n1156));
  NAND4_X1  g730(.A1(new_n949), .A2(new_n880), .A3(new_n694), .A4(new_n1156), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


