//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n209), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT65), .Z(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  AND2_X1   g0024(.A1(KEYINPUT67), .A2(G77), .ZN(new_n225));
  NOR2_X1   g0025(.A1(KEYINPUT67), .A2(G77), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n223), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n229), .B(new_n230), .C1(new_n201), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n206), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n221), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n211), .A2(new_n213), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n258), .A2(new_n216), .A3(G1), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR3_X1   g0063(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G150), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n261), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT70), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OR3_X1    g0070(.A1(new_n269), .A2(new_n201), .A3(KEYINPUT8), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n216), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n267), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n211), .A2(new_n213), .A3(new_n252), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n257), .B1(G50), .B2(new_n260), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  XOR2_X1   g0079(.A(new_n279), .B(KEYINPUT9), .Z(new_n280));
  OAI21_X1  g0080(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  INV_X1    g0087(.A(G226), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n214), .A2(new_n285), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G222), .A2(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G223), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n227), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n293), .B(new_n302), .C1(new_n303), .C2(new_n298), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n289), .A2(new_n290), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n291), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n306), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n280), .B2(new_n309), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n279), .C1(G179), .C2(new_n306), .ZN(new_n315));
  INV_X1    g0115(.A(new_n287), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n283), .B1(new_n316), .B2(G244), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n298), .A2(G232), .A3(new_n300), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT72), .B(G107), .Z(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n298), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n300), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n320), .B1(G238), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n317), .B1(new_n325), .B2(new_n292), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G179), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT74), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT71), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(new_n216), .A3(new_n295), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n262), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n268), .B1(new_n331), .B2(KEYINPUT73), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(KEYINPUT73), .B2(new_n331), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT15), .B(G87), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n333), .B1(new_n216), .B2(new_n227), .C1(new_n274), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n277), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n256), .A2(G77), .B1(new_n227), .B2(new_n259), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(new_n337), .B1(new_n326), .B2(new_n313), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n326), .A2(new_n308), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n326), .A2(G200), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n340), .A2(new_n336), .A3(new_n337), .A4(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n312), .A2(new_n315), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n253), .A2(new_n202), .A3(G13), .A4(G20), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT76), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(new_n346), .C1(new_n202), .C2(new_n255), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT12), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n344), .B(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n255), .A2(new_n202), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT76), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G50), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n330), .B2(new_n262), .ZN(new_n354));
  INV_X1    g0154(.A(G77), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n274), .A2(new_n355), .B1(new_n216), .B2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n277), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT11), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT11), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n277), .C1(new_n354), .C2(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT77), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(G226), .B(new_n300), .C1(new_n321), .C2(new_n322), .ZN(new_n367));
  OAI211_X1 g0167(.A(G232), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n367), .A2(new_n368), .A3(new_n372), .A4(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n373), .A3(new_n293), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT13), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n283), .B1(new_n316), .B2(G238), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n374), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g0179(.A(G200), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n374), .A2(new_n376), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(G190), .A3(new_n377), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n366), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n366), .A2(new_n380), .A3(KEYINPUT78), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n272), .B1(new_n253), .B2(G20), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n277), .A2(new_n259), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n390), .A2(new_n391), .B1(new_n259), .B2(new_n272), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n216), .B1(new_n203), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT80), .B1(new_n331), .B2(G159), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT80), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n330), .C2(new_n262), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n323), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n296), .A2(new_n216), .A3(new_n297), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n403), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n401), .B1(new_n408), .B2(G68), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n410));
  NAND2_X1  g0210(.A1(new_n403), .A2(new_n405), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n202), .B1(new_n411), .B2(new_n402), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n409), .A2(KEYINPUT16), .B1(new_n413), .B2(KEYINPUT82), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n398), .B1(new_n265), .B2(new_n399), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n331), .A2(KEYINPUT80), .A3(G159), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n395), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n412), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT82), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n278), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n393), .B1(new_n414), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n284), .B1(new_n287), .B2(new_n231), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n288), .A2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G223), .B2(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G87), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n426), .A2(new_n323), .B1(new_n295), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n428), .B2(new_n293), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n313), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(G179), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT18), .B1(new_n423), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n402), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n418), .B(KEYINPUT16), .C1(new_n436), .C2(new_n202), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n420), .B2(new_n421), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n277), .B1(new_n413), .B2(KEYINPUT82), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n392), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n431), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n378), .A2(new_n379), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT14), .B1(new_n446), .B2(new_n313), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT14), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(G169), .C1(new_n378), .C2(new_n379), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(G179), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n366), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n429), .A2(new_n308), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(G200), .B2(new_n429), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n392), .B(new_n455), .C1(new_n438), .C2(new_n439), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n414), .A2(new_n422), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(KEYINPUT17), .A3(new_n392), .A4(new_n455), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n445), .A2(new_n453), .A3(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n343), .A2(new_n389), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G244), .B(new_n300), .C1(new_n321), .C2(new_n322), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n298), .A2(KEYINPUT4), .A3(G244), .A4(new_n300), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n298), .A2(G250), .A3(G1698), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n293), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n472), .A2(G274), .A3(new_n286), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n474), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n476), .A2(G257), .A3(new_n286), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n471), .A2(new_n308), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n475), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n480), .B(new_n477), .C1(new_n470), .C2(new_n293), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(G200), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n483), .A2(new_n484), .A3(G107), .ZN(new_n485));
  XNOR2_X1  g0285(.A(G97), .B(G107), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n487), .A2(new_n216), .B1(new_n355), .B2(new_n265), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n319), .B1(new_n411), .B2(new_n402), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n277), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n260), .A2(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n295), .A2(G1), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n277), .A2(new_n259), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(KEYINPUT83), .A3(new_n494), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n482), .A2(KEYINPUT84), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n477), .B1(new_n470), .B2(new_n293), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n475), .ZN(new_n501));
  INV_X1    g0301(.A(G179), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n313), .B1(new_n500), .B2(new_n475), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n495), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n490), .A2(KEYINPUT83), .A3(new_n494), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT83), .B1(new_n490), .B2(new_n494), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT84), .B1(new_n509), .B2(new_n482), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(G20), .B1(G33), .B2(G283), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n295), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n512), .A2(new_n513), .B1(G20), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT90), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n277), .B1(new_n516), .B2(KEYINPUT20), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n516), .B2(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n493), .A2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n259), .A2(new_n514), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT20), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n515), .A2(new_n277), .A3(KEYINPUT90), .A4(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(new_n300), .C1(new_n321), .C2(new_n322), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT88), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT89), .B(G303), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n324), .A2(G264), .B1(new_n323), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n292), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n476), .A2(G270), .A3(new_n286), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n475), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n523), .B(G169), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n529), .A2(new_n502), .A3(new_n531), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n523), .ZN(new_n535));
  INV_X1    g0335(.A(new_n531), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n526), .A2(new_n528), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n292), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT21), .A3(G169), .A4(new_n523), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n216), .B(G87), .C1(new_n321), .C2(new_n322), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT22), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n216), .A2(KEYINPUT23), .A3(G107), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT72), .B(G107), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(KEYINPUT23), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT91), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n295), .A2(new_n514), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n216), .B1(new_n547), .B2(KEYINPUT23), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT24), .B(new_n542), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n278), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n493), .A2(G107), .ZN(new_n555));
  INV_X1    g0355(.A(G107), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n259), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT25), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT92), .ZN(new_n559));
  OR3_X1    g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n555), .B2(new_n558), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n551), .A2(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n476), .A2(G264), .A3(new_n286), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n475), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n298), .A2(G257), .A3(G1698), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n298), .A2(G250), .A3(new_n300), .ZN(new_n566));
  INV_X1    g0366(.A(G294), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n566), .C1(new_n295), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n564), .B1(new_n293), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n502), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n569), .B2(G169), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n540), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n538), .A2(G200), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n529), .A2(new_n531), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  INV_X1    g0376(.A(new_n523), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n554), .A2(new_n551), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n560), .A2(new_n561), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n569), .A2(G190), .ZN(new_n582));
  INV_X1    g0382(.A(G200), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(new_n569), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n578), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n298), .A2(G244), .A3(G1698), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n298), .A2(G238), .A3(new_n300), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n293), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n253), .A2(G45), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n286), .A2(G250), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n474), .B2(G274), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n286), .A2(new_n593), .A3(G250), .A4(new_n591), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT86), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n590), .B(new_n502), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G87), .A2(G97), .ZN(new_n601));
  NAND3_X1  g0401(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n319), .A2(new_n601), .B1(new_n216), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n216), .B(G68), .C1(new_n321), .C2(new_n322), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n274), .B2(new_n484), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n277), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n334), .A2(new_n259), .ZN(new_n609));
  INV_X1    g0409(.A(new_n334), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n493), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n595), .A2(new_n596), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT86), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n615), .B1(new_n293), .B2(new_n589), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n600), .B(new_n612), .C1(new_n616), .C2(G169), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n590), .B(G190), .C1(new_n598), .C2(new_n599), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n493), .A2(G87), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n608), .A2(new_n609), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(G200), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n618), .B1(new_n622), .B2(KEYINPUT87), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT87), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n624), .B(new_n620), .C1(G200), .C2(new_n621), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n617), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n585), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n463), .A2(new_n511), .A3(new_n573), .A4(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n384), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n453), .B1(new_n629), .B2(new_n339), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n461), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n312), .B1(new_n631), .B2(new_n444), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n315), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n608), .A2(new_n609), .A3(new_n619), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n635), .B(new_n618), .C1(new_n616), .C2(new_n583), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n617), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT93), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT93), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n617), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n535), .B(new_n539), .C1(new_n562), .C2(new_n571), .ZN(new_n642));
  INV_X1    g0442(.A(new_n584), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n562), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n510), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n499), .A3(new_n505), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT94), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n638), .A2(new_n640), .B1(new_n562), .B2(new_n643), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT94), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n511), .A2(new_n649), .A3(new_n650), .A4(new_n642), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n501), .A2(G169), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n481), .A2(G179), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n654), .A2(new_n655), .B1(new_n497), .B2(new_n498), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n641), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n495), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n655), .B2(new_n654), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n659), .B(new_n617), .C1(new_n623), .C2(new_n625), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n657), .A2(new_n617), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n463), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n634), .A2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n253), .A2(new_n216), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n577), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n540), .B(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(new_n578), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n644), .B1(new_n562), .B2(new_n672), .ZN(new_n677));
  INV_X1    g0477(.A(new_n572), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n572), .A2(new_n672), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n540), .A2(new_n672), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n680), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n207), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G1), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n319), .A2(new_n514), .A3(new_n601), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n218), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT98), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n511), .A2(new_n649), .A3(new_n642), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT96), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n660), .A2(new_n698), .A3(new_n653), .ZN(new_n699));
  INV_X1    g0499(.A(new_n640), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n639), .B1(new_n617), .B2(new_n636), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT26), .B(new_n656), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n660), .B2(new_n653), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n697), .B(new_n617), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT97), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n705), .A2(new_n706), .A3(new_n672), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n705), .B2(new_n672), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n696), .B(KEYINPUT29), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n672), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(new_n706), .A3(new_n672), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n671), .B1(new_n652), .B2(new_n662), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT98), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n709), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n627), .A2(new_n511), .A3(new_n573), .A4(new_n672), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n575), .A2(G179), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n616), .A2(new_n569), .A3(new_n500), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n723), .A2(new_n724), .A3(new_n722), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(KEYINPUT95), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n569), .A2(G179), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n538), .A2(new_n729), .A3(new_n501), .A4(new_n621), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n725), .B2(KEYINPUT95), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n671), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n726), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n725), .A3(new_n730), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n719), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n718), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n695), .B1(new_n740), .B2(G1), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT99), .Z(G364));
  NOR2_X1   g0542(.A1(new_n258), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n253), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n690), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n676), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n675), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n748), .B1(new_n719), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n216), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT100), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n215), .B1(G20), .B2(new_n313), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n753), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT101), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n689), .A2(new_n323), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G355), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G116), .B2(new_n207), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n247), .A2(new_n473), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n298), .B(new_n689), .C1(new_n219), .C2(new_n473), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n746), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT102), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n216), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G159), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT32), .Z(new_n773));
  NOR2_X1   g0573(.A1(new_n216), .A2(new_n308), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n502), .A2(new_n583), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n583), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n777), .A2(G50), .B1(new_n780), .B2(G107), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n502), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n769), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n227), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n774), .A2(new_n778), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n298), .B1(new_n785), .B2(new_n427), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n782), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n775), .A2(new_n769), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n201), .A2(new_n787), .B1(new_n788), .B2(new_n202), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n784), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(G20), .B1(new_n768), .B2(new_n308), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G97), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n773), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT103), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n788), .B1(new_n795), .B2(KEYINPUT103), .ZN(new_n797));
  INV_X1    g0597(.A(new_n787), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(new_n797), .B1(G322), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT104), .Z(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n785), .A2(new_n801), .B1(new_n783), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G326), .B2(new_n777), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n791), .A2(G294), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n771), .A2(G329), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n298), .B1(new_n780), .B2(G283), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n793), .B1(new_n800), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n766), .B1(new_n809), .B2(new_n756), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n750), .B1(new_n755), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n339), .A2(new_n671), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n336), .A2(new_n337), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n671), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n342), .A2(new_n815), .B1(new_n328), .B2(new_n338), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n715), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n746), .B1(new_n818), .B2(new_n738), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n738), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n756), .A2(new_n751), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G77), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n776), .A2(new_n801), .B1(new_n788), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n785), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G107), .B2(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n787), .A2(new_n567), .B1(new_n783), .B2(new_n514), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n779), .A2(new_n427), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n828), .A2(new_n298), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n771), .A2(G311), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n830), .A3(new_n792), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n783), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G143), .A2(new_n798), .B1(new_n833), .B2(G159), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n835), .B2(new_n776), .C1(new_n266), .C2(new_n788), .ZN(new_n836));
  XOR2_X1   g0636(.A(KEYINPUT105), .B(KEYINPUT34), .Z(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n298), .B1(new_n785), .B2(new_n353), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G68), .B2(new_n780), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  INV_X1    g0641(.A(new_n771), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n838), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n791), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n836), .A2(new_n837), .B1(new_n201), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n832), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n747), .B(new_n823), .C1(new_n846), .C2(new_n756), .ZN(new_n847));
  INV_X1    g0647(.A(new_n751), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n817), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n820), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  INV_X1    g0651(.A(new_n487), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(G116), .A3(new_n217), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  NAND3_X1  g0656(.A1(new_n219), .A2(new_n303), .A3(new_n394), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n353), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n253), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n813), .B(KEYINPUT106), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n715), .B2(new_n817), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n452), .A2(new_n671), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n453), .A2(new_n384), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT107), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n451), .B1(new_n386), .B2(new_n387), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n864), .B(new_n865), .C1(new_n863), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n451), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n863), .B1(new_n388), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n863), .A2(new_n384), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n452), .B2(new_n451), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT107), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n432), .A2(new_n443), .A3(new_n458), .A4(new_n460), .ZN(new_n875));
  INV_X1    g0675(.A(new_n437), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n277), .B1(new_n409), .B2(new_n415), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT108), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n418), .B1(new_n436), .B2(new_n202), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n278), .B1(new_n880), .B2(new_n410), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT108), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n393), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n669), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n875), .A2(KEYINPUT109), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT109), .B1(new_n875), .B2(new_n884), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  INV_X1    g0687(.A(new_n456), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n437), .B1(new_n881), .B2(KEYINPUT108), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n877), .A2(new_n878), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n392), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n669), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n441), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n440), .A2(new_n441), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n440), .A2(new_n892), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(new_n456), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n885), .A2(new_n886), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n456), .B1(new_n883), .B2(new_n669), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n883), .A2(new_n431), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n907), .B(KEYINPUT38), .C1(new_n886), .C2(new_n885), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n874), .A2(new_n909), .B1(new_n444), .B2(new_n669), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n451), .A2(new_n452), .A3(new_n672), .ZN(new_n912));
  INV_X1    g0712(.A(new_n908), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n875), .A2(new_n884), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT109), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n875), .A2(KEYINPUT109), .A3(new_n884), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n918), .B2(new_n907), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT39), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT110), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n898), .B(new_n887), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n897), .B1(new_n445), .B2(new_n461), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n901), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n908), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n920), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n902), .B2(new_n908), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n908), .A2(new_n922), .A3(new_n925), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT110), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n912), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n911), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n633), .B1(new_n717), .B2(new_n463), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n731), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n672), .B1(new_n935), .B2(new_n727), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n720), .B2(KEYINPUT31), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(KEYINPUT31), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n817), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n873), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n909), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n908), .B2(new_n925), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n941), .A2(new_n942), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n937), .A2(new_n938), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n944), .A2(new_n463), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n463), .B2(new_n945), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n946), .A2(new_n947), .A3(new_n719), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n934), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n253), .B2(new_n743), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n934), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n860), .B1(new_n950), .B2(new_n951), .ZN(G367));
  INV_X1    g0752(.A(new_n685), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n681), .A2(new_n684), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n676), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n718), .A2(new_n738), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT112), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n953), .A2(new_n680), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n511), .B1(new_n509), .B2(new_n672), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n656), .A2(new_n671), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n961), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT45), .B1(new_n687), .B2(new_n964), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT44), .B1(new_n961), .B2(new_n965), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT44), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n687), .A2(new_n970), .A3(new_n964), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n967), .A2(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n683), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n959), .A2(new_n960), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n682), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT112), .B1(new_n975), .B2(new_n958), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n739), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n690), .B(KEYINPUT41), .Z(new_n978));
  OAI21_X1  g0778(.A(new_n744), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n682), .A2(new_n964), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT111), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n641), .B1(new_n635), .B2(new_n672), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n617), .A2(new_n635), .A3(new_n672), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n685), .A2(new_n964), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n964), .A2(new_n572), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n671), .B1(new_n988), .B2(new_n505), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n985), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n981), .B(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n979), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n689), .A2(new_n298), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n243), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n207), .B2(new_n334), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n746), .B1(new_n759), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT46), .B1(new_n826), .B2(G116), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT113), .Z(new_n1000));
  NAND3_X1  g0800(.A1(new_n826), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(new_n323), .C1(new_n824), .C2(new_n783), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n527), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1003), .A2(new_n787), .B1(new_n788), .B2(new_n567), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n780), .A2(G97), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n802), .B2(new_n776), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT114), .B(G317), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n771), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n791), .A2(new_n544), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1000), .A2(new_n1007), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n842), .A2(new_n835), .B1(new_n201), .B2(new_n785), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n266), .A2(new_n787), .B1(new_n788), .B2(new_n399), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n227), .A2(new_n779), .B1(new_n783), .B2(new_n353), .ZN(new_n1016));
  INV_X1    g0816(.A(G143), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n298), .B1(new_n776), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1014), .B(new_n1019), .C1(new_n202), .C2(new_n844), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1011), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n998), .B1(new_n1023), .B2(new_n756), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n984), .B2(new_n753), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n994), .A2(new_n1025), .ZN(G387));
  NAND3_X1  g0826(.A1(new_n958), .A2(KEYINPUT116), .A3(new_n690), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n958), .A2(new_n690), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT116), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1027), .B(new_n1030), .C1(new_n740), .C2(new_n957), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n323), .B1(new_n779), .B2(new_n514), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n788), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n777), .A2(G322), .B1(new_n1033), .B2(G311), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n798), .A2(new_n1008), .B1(new_n833), .B2(new_n527), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n824), .B2(new_n844), .C1(new_n567), .C2(new_n785), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT49), .Z(new_n1039));
  AOI211_X1 g0839(.A(new_n1032), .B(new_n1039), .C1(G326), .C2(new_n771), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G159), .A2(new_n777), .B1(new_n826), .B2(new_n303), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G50), .A2(new_n798), .B1(new_n833), .B2(G68), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1041), .A2(new_n1042), .A3(new_n298), .A4(new_n1005), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n842), .A2(new_n266), .B1(new_n272), .B2(new_n788), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n844), .A2(new_n334), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n756), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n240), .A2(G45), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(new_n995), .B1(new_n693), .B2(new_n760), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n268), .A2(G50), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT50), .Z(new_n1051));
  OAI21_X1  g0851(.A(new_n473), .B1(new_n202), .B2(new_n355), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1051), .A2(new_n693), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n556), .B2(new_n689), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1047), .B(new_n746), .C1(new_n759), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n681), .B2(new_n754), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n957), .B2(new_n745), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1031), .A2(new_n1058), .ZN(G393));
  NAND2_X1  g0859(.A1(new_n965), .A2(new_n754), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT117), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n250), .A2(new_n995), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n484), .B2(new_n207), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n746), .B1(new_n759), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G317), .A2(new_n777), .B1(new_n798), .B2(G311), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT52), .Z(new_n1066));
  OAI22_X1  g0866(.A1(new_n1003), .A2(new_n788), .B1(new_n783), .B2(new_n567), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n298), .B(new_n1067), .C1(G107), .C2(new_n780), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(new_n514), .C2(new_n844), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n771), .A2(G322), .B1(G283), .B2(new_n826), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT118), .Z(new_n1071));
  NOR2_X1   g0871(.A1(new_n844), .A2(new_n355), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G50), .A2(new_n1033), .B1(new_n826), .B2(G68), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n268), .B2(new_n783), .ZN(new_n1074));
  OR4_X1    g0874(.A1(new_n323), .A2(new_n1072), .A3(new_n1074), .A4(new_n829), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G150), .A2(new_n777), .B1(new_n798), .B2(G159), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(KEYINPUT51), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n1017), .C2(new_n842), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1069), .A2(new_n1071), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1064), .B1(new_n1080), .B2(new_n756), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1061), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n975), .B2(new_n744), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n974), .A2(new_n976), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n691), .B1(new_n975), .B2(new_n958), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(G390));
  OAI21_X1  g0887(.A(new_n912), .B1(new_n862), .B2(new_n873), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n927), .A2(new_n930), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n912), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n908), .B2(new_n925), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n712), .A2(new_n713), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n861), .B1(new_n1092), .B2(new_n817), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1093), .B2(new_n873), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n939), .A2(new_n873), .A3(new_n719), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n945), .A2(new_n463), .A3(G330), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n933), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n736), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n817), .C1(new_n937), .C2(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(new_n873), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1089), .A2(new_n1094), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n862), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1101), .A2(new_n873), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n1096), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n817), .B1(new_n707), .B2(new_n708), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n861), .ZN(new_n1108));
  OAI211_X1 g0908(.A(G330), .B(new_n817), .C1(new_n937), .C2(new_n938), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n873), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1102), .A2(new_n1107), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1097), .A2(new_n1099), .A3(new_n1103), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n717), .A2(new_n463), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1112), .A2(new_n1114), .A3(new_n634), .A4(new_n1098), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1089), .A2(new_n1094), .A3(new_n1102), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1096), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1115), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1113), .A2(new_n1119), .A3(new_n690), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1097), .A2(new_n745), .A3(new_n1103), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n746), .B1(new_n822), .B2(new_n273), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G128), .A2(new_n777), .B1(new_n798), .B2(G132), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT119), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n399), .B2(new_n844), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n785), .A2(new_n266), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n771), .A2(G125), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n323), .B1(new_n780), .B2(G50), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G137), .A2(new_n1033), .B1(new_n833), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n202), .A2(new_n779), .B1(new_n783), .B2(new_n484), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n298), .B(new_n1134), .C1(G87), .C2(new_n826), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n776), .A2(new_n824), .B1(new_n787), .B2(new_n514), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n544), .B2(new_n1033), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n567), .C2(new_n842), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1125), .A2(new_n1133), .B1(new_n1138), .B2(new_n1072), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1122), .B1(new_n1139), .B2(new_n756), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT110), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n921), .B1(new_n920), .B2(new_n926), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1140), .B1(new_n1144), .B2(new_n848), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1120), .A2(new_n1121), .A3(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n941), .A2(new_n942), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n279), .A2(new_n892), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n312), .A2(new_n315), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n312), .B2(new_n315), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n943), .A2(new_n940), .ZN(new_n1157));
  AND4_X1   g0957(.A1(G330), .A2(new_n1147), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n944), .B2(G330), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1158), .A2(new_n1159), .B1(new_n931), .B2(new_n911), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1147), .A2(G330), .A3(new_n1157), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1156), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1090), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n944), .A2(G330), .A3(new_n1156), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n910), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1116), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n933), .A2(new_n1098), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(KEYINPUT57), .B(new_n1167), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n690), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1162), .A2(new_n751), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n746), .B1(new_n822), .B2(G50), .ZN(new_n1176));
  INV_X1    g0976(.A(G41), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G50), .B1(new_n297), .B2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n484), .A2(new_n788), .B1(new_n787), .B2(new_n556), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n777), .A2(G116), .B1(new_n833), .B2(new_n610), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n201), .B2(new_n779), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G68), .C2(new_n791), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1177), .B(new_n323), .C1(new_n785), .C2(new_n227), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT120), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n824), .C2(new_n842), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1178), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n788), .A2(new_n841), .B1(new_n783), .B2(new_n835), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT121), .Z(new_n1189));
  AOI22_X1  g0989(.A1(G125), .A2(new_n777), .B1(new_n798), .B2(G128), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT122), .B1(new_n785), .B2(new_n1130), .ZN(new_n1191));
  OR3_X1    g0991(.A1(new_n785), .A2(new_n1130), .A3(KEYINPUT122), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1189), .B(new_n1193), .C1(new_n266), .C2(new_n844), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n295), .B(new_n1177), .C1(new_n779), .C2(new_n399), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n771), .B2(G124), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1176), .B1(new_n1200), .B2(new_n756), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1167), .A2(new_n745), .B1(new_n1175), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1174), .A2(new_n1202), .ZN(G375));
  NAND3_X1  g1003(.A1(new_n1169), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n978), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1115), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n873), .A2(new_n751), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n746), .B1(new_n822), .B2(G68), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n776), .A2(new_n841), .B1(new_n788), .B2(new_n1130), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n323), .B(new_n1209), .C1(G58), .C2(new_n780), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n791), .A2(G50), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n771), .A2(G128), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n787), .A2(new_n835), .B1(new_n783), .B2(new_n266), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G159), .B2(new_n826), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n319), .A2(new_n783), .B1(new_n779), .B2(new_n355), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n298), .B(new_n1216), .C1(G294), .C2(new_n777), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n514), .A2(new_n788), .B1(new_n787), .B2(new_n824), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G97), .B2(new_n826), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(new_n801), .C2(new_n842), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1215), .B1(new_n1220), .B2(new_n1045), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT123), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n757), .B1(new_n1221), .B2(KEYINPUT123), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1208), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1112), .A2(new_n745), .B1(new_n1207), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1225), .ZN(G381));
  AND2_X1   g1026(.A1(new_n1174), .A2(new_n1202), .ZN(new_n1227));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1031), .A2(new_n811), .A3(new_n1058), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1229), .A2(new_n1231), .A3(G387), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT124), .Z(G407));
  INV_X1    g1033(.A(G213), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1229), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(G343), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT125), .Z(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G407), .A2(new_n1238), .ZN(G409));
  NAND2_X1  g1039(.A1(new_n1115), .A2(KEYINPUT60), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n690), .B1(new_n1204), .B2(new_n1240), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1204), .A2(new_n1240), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1225), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(new_n850), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n850), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT61), .B1(new_n1246), .B2(KEYINPUT62), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1173), .A2(new_n690), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1113), .A2(new_n1099), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1167), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G378), .B(new_n1202), .C1(new_n1248), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT126), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT126), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1174), .A2(new_n1253), .A3(G378), .A4(new_n1202), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1202), .B1(new_n1170), .B2(new_n978), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1228), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1237), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1236), .A2(G2897), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1244), .A2(new_n1245), .A3(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1244), .A2(new_n1245), .B1(G2897), .B2(new_n1237), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1260), .A2(new_n1261), .A3(KEYINPUT62), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1247), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1252), .A2(new_n1254), .B1(new_n1228), .B2(new_n1256), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1264), .A2(KEYINPUT62), .A3(new_n1236), .A4(new_n1246), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n994), .A2(new_n1025), .A3(G390), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G390), .B1(new_n994), .B2(new_n1025), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1230), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n811), .B1(new_n1031), .B2(new_n1058), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1268), .A2(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1269), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1267), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1264), .A2(new_n1236), .B1(new_n1261), .B2(new_n1260), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1246), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1236), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1277), .A2(KEYINPUT63), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(KEYINPUT61), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1278), .A2(KEYINPUT63), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1258), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1266), .A2(new_n1276), .B1(new_n1280), .B2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1228), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1255), .A2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1276), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(new_n1281), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1287), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1276), .A2(new_n1289), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1281), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(KEYINPUT127), .A4(new_n1278), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(G402));
endmodule


