//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n466), .B2(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n467), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n471), .A2(new_n476), .A3(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n470), .A2(new_n465), .A3(G2105), .A4(new_n467), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n470), .A2(new_n465), .A3(new_n469), .A4(new_n467), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(new_n486), .B2(G136), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n470), .A2(new_n465), .A3(new_n467), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n472), .A2(new_n467), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n488), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n469), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT67), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(new_n496), .B2(new_n497), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n470), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XOR2_X1   g079(.A(KEYINPUT6), .B(G651), .Z(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT68), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n508), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(G50), .A2(new_n517), .B1(new_n520), .B2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XNOR2_X1  g098(.A(KEYINPUT69), .B(G51), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n517), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n510), .A2(G63), .ZN(new_n528));
  AND3_X1   g103(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(G651), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n509), .A2(G89), .A3(new_n513), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT70), .ZN(new_n535));
  INV_X1    g110(.A(G77), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI221_X1 g112(.A(KEYINPUT70), .B1(new_n536), .B2(new_n516), .C1(new_n508), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(G651), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n514), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n517), .A2(G52), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n514), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n508), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(G43), .A2(new_n517), .B1(new_n547), .B2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n511), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n511), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G651), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n509), .A2(G91), .A3(new_n513), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(new_n531), .B2(new_n532), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g146(.A1(new_n531), .A2(new_n569), .A3(new_n532), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(G286));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n565), .B1(new_n508), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n517), .B2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n509), .A2(new_n513), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(G288));
  OAI21_X1  g154(.A(G61), .B1(new_n506), .B2(new_n507), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n565), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(KEYINPUT74), .A2(new_n582), .B1(new_n517), .B2(G48), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n582), .A2(KEYINPUT74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n509), .A2(G86), .A3(new_n513), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n514), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(G651), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n565), .B1(new_n595), .B2(new_n558), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n577), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  MUX2_X1   g185(.A(new_n607), .B(new_n609), .S(new_n610), .Z(G297));
  MUX2_X1   g186(.A(new_n607), .B(new_n609), .S(new_n610), .Z(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n604), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n492), .A2(new_n477), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n623), .A2(new_n624), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n624), .B2(new_n623), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n480), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n486), .B2(G135), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n622), .A2(new_n632), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT79), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n652), .A2(new_n655), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n652), .A2(new_n655), .A3(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT83), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT84), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT85), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  INV_X1    g267(.A(G288), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(new_n688), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n688), .B2(G23), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(G6), .A2(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G305), .B2(new_n688), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n695), .A2(new_n696), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n697), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n692), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT34), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n692), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  INV_X1    g286(.A(G95), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n712), .A2(new_n469), .A3(KEYINPUT86), .ZN(new_n713));
  AOI21_X1  g288(.A(KEYINPUT86), .B1(new_n712), .B2(new_n469), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G107), .B2(new_n469), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G119), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n480), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n486), .A2(G131), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n711), .B1(new_n719), .B2(new_n710), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT87), .B(G1986), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n707), .A2(new_n709), .A3(new_n722), .A4(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(new_n469), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT91), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT25), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n486), .B2(G139), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n710), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n710), .B2(G33), .ZN(new_n738));
  INV_X1    g313(.A(G2072), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT24), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(KEYINPUT24), .ZN(new_n742));
  AOI22_X1  g317(.A1(G160), .A2(G29), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n738), .A2(new_n739), .B1(G2084), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT27), .B(G1996), .Z(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT26), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(new_n477), .B2(G105), .ZN(new_n750));
  INV_X1    g325(.A(G129), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n480), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G141), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n485), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n752), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n760), .B(new_n761), .C1(G29), .C2(G32), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n744), .B1(new_n739), .B2(new_n738), .C1(new_n745), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G19), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n550), .B2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G1341), .Z(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G168), .A2(new_n688), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n688), .B2(G21), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n768), .B1(new_n769), .B2(new_n771), .C1(G2084), .C2(new_n743), .ZN(new_n772));
  NOR2_X1   g347(.A1(G5), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G171), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT96), .B(G1961), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n604), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT89), .B(G1348), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n771), .A2(new_n769), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT95), .B(G28), .Z(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n783), .B(new_n788), .C1(new_n710), .C2(new_n631), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n688), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT23), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n608), .B2(new_n688), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n710), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT28), .ZN(new_n796));
  INV_X1    g371(.A(G104), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n797), .A2(new_n469), .A3(KEYINPUT90), .ZN(new_n798));
  AOI21_X1  g373(.A(KEYINPUT90), .B1(new_n797), .B2(new_n469), .ZN(new_n799));
  OAI221_X1 g374(.A(G2104), .B1(G116), .B2(new_n469), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G128), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n480), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n486), .A2(G140), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n796), .B1(new_n804), .B2(new_n710), .ZN(new_n805));
  INV_X1    g380(.A(G2067), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n794), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n772), .A2(new_n782), .A3(new_n789), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G29), .A2(G35), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G162), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT29), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2090), .ZN(new_n813));
  NOR2_X1   g388(.A1(G27), .A2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G164), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2078), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n813), .B(new_n817), .C1(new_n745), .C2(new_n763), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n765), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n728), .A2(new_n819), .ZN(G311));
  INV_X1    g395(.A(G311), .ZN(G150));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n549), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n565), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT98), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n514), .A2(G93), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT99), .B(G55), .Z(new_n828));
  AOI22_X1  g403(.A1(new_n825), .A2(KEYINPUT98), .B1(new_n517), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n544), .A2(KEYINPUT100), .A3(new_n548), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n823), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(new_n822), .A3(new_n549), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n600), .A2(new_n603), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n596), .B(new_n597), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n613), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n836), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n833), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n495), .A2(new_n848), .A3(new_n501), .A4(new_n502), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT67), .ZN(new_n850));
  INV_X1    g425(.A(new_n497), .ZN(new_n851));
  INV_X1    g426(.A(G114), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G2105), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G126), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n854), .A2(new_n498), .B1(new_n480), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT101), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n486), .A2(G142), .ZN(new_n860));
  INV_X1    g435(.A(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n469), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n860), .B1(new_n861), .B2(new_n480), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n620), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n759), .A2(new_n804), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n758), .A2(new_n803), .A3(new_n802), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n719), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n867), .A2(new_n868), .A3(new_n719), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n865), .A3(new_n869), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n859), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n874), .A3(new_n859), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(new_n736), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n735), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n630), .B(G160), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G162), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n878), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G395));
  NAND2_X1  g464(.A1(new_n832), .A2(new_n834), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n615), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n604), .B2(G299), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n839), .A2(KEYINPUT103), .A3(new_n608), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n837), .A2(new_n838), .A3(G299), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT102), .B1(new_n604), .B2(G299), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n893), .B(new_n894), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n895), .B(new_n896), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n893), .A4(new_n894), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n906), .B2(new_n891), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n908));
  XNOR2_X1  g483(.A(G290), .B(G305), .ZN(new_n909));
  XNOR2_X1  g484(.A(G303), .B(new_n693), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n908), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g491(.A(new_n915), .B1(G868), .B2(new_n830), .ZN(G331));
  NAND2_X1  g492(.A1(G168), .A2(KEYINPUT73), .ZN(new_n918));
  AOI21_X1  g493(.A(G301), .B1(new_n918), .B2(new_n570), .ZN(new_n919));
  NOR2_X1   g494(.A1(G171), .A2(G168), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n890), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(G171), .B1(new_n571), .B2(new_n572), .ZN(new_n922));
  INV_X1    g497(.A(G168), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G301), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n922), .A2(new_n832), .A3(new_n834), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n902), .A2(new_n905), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n911), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n919), .A2(new_n920), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n835), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(KEYINPUT105), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n899), .A4(new_n921), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n928), .B1(new_n927), .B2(new_n933), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n899), .A2(new_n921), .A3(KEYINPUT106), .A4(new_n925), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n899), .A2(new_n921), .A3(new_n925), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n931), .A2(new_n932), .A3(new_n921), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n902), .A2(new_n905), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n942), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n936), .B1(new_n911), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n940), .B(KEYINPUT44), .C1(new_n941), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n911), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(new_n935), .A3(new_n937), .A4(new_n934), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT107), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n957), .B(KEYINPUT44), .C1(new_n952), .C2(new_n953), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n956), .B2(new_n958), .ZN(G397));
  INV_X1    g534(.A(new_n859), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT108), .B(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND4_X1   g537(.A1(G40), .A2(new_n471), .A3(new_n476), .A4(new_n478), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT110), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AND4_X1   g542(.A1(KEYINPUT110), .A2(new_n962), .A3(new_n966), .A4(new_n963), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n759), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n804), .B(G2067), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n966), .B2(new_n759), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n721), .A3(new_n719), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n804), .A2(new_n806), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n972), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n719), .B(new_n721), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n964), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n965), .A2(G1986), .A3(G290), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT48), .Z(new_n980));
  AND2_X1   g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n965), .B1(new_n759), .B2(new_n970), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n967), .A2(new_n983), .A3(new_n968), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n967), .B2(new_n968), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n975), .B(new_n981), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n963), .A2(new_n991), .A3(new_n503), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n576), .B(G1976), .C1(new_n577), .C2(new_n578), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(G8), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT52), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(new_n992), .A3(G8), .A4(new_n993), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n992), .A2(G8), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n583), .A2(new_n584), .A3(new_n1002), .A4(new_n585), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n1005), .B2(KEYINPUT49), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n999), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n471), .A2(new_n476), .A3(G40), .A4(new_n478), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n991), .B1(new_n856), .B2(new_n857), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n849), .A2(new_n858), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G2078), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n503), .A2(new_n1019), .A3(new_n991), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n963), .ZN(new_n1022));
  INV_X1    g597(.A(G1961), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1017), .A2(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1018), .A2(G2078), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1013), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G301), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1022), .A2(G2090), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1030));
  OAI21_X1  g605(.A(G8), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n515), .B2(new_n521), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(G8), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1009), .A2(new_n1028), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G168), .A2(new_n1032), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1013), .A2(new_n1026), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n769), .ZN(new_n1046));
  INV_X1    g621(.A(G2084), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1020), .A2(new_n1021), .A3(new_n1047), .A4(new_n963), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1044), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT51), .B1(new_n1043), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1032), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(new_n1043), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1048), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1966), .B1(new_n1013), .B2(new_n1026), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n1044), .A3(new_n1051), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1049), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1041), .B1(new_n1042), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1049), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1053), .A2(new_n1052), .A3(new_n1043), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1051), .B1(new_n1057), .B2(new_n1044), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1059), .B2(new_n1042), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1060), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT126), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1060), .A2(new_n1065), .A3(new_n1067), .A4(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(new_n1003), .B(KEYINPUT113), .Z(new_n1072));
  NAND2_X1  g647(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G288), .A2(G1976), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT114), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1009), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1076), .A2(new_n1000), .B1(new_n1077), .B2(new_n1040), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1037), .B1(new_n1031), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1079), .B2(new_n1031), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1057), .A2(new_n1082), .A3(G286), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1081), .A2(new_n1040), .A3(new_n1009), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1057), .A2(G286), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1009), .A2(new_n1085), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1082), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1078), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1069), .A2(new_n1071), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1015), .A2(new_n963), .A3(new_n1025), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n962), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1024), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT124), .B1(new_n1092), .B2(G171), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1028), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G301), .A4(new_n1024), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1092), .A2(G171), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1024), .A2(G301), .A3(new_n1027), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(KEYINPUT54), .A3(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1009), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1099), .A2(new_n1102), .A3(new_n1103), .A4(new_n1064), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1013), .A2(new_n1015), .A3(new_n966), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1013), .A2(new_n1015), .A3(new_n1110), .A4(new_n966), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n992), .A2(KEYINPUT119), .A3(new_n1112), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n550), .B(new_n1106), .C1(new_n1109), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1108), .A2(new_n1111), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1106), .B1(new_n1120), .B2(new_n550), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n608), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1022), .A2(new_n793), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1013), .A2(new_n1015), .A3(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1123), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1125), .A2(new_n1138), .A3(new_n1126), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT61), .B(new_n1135), .C1(new_n1136), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n1122), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n550), .B1(new_n1109), .B2(new_n1117), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1105), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1118), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n1134), .A4(new_n1141), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n963), .A2(new_n991), .A3(new_n806), .A4(new_n503), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT116), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(G1348), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1022), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1149), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1154), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n604), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n839), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1143), .A2(new_n1148), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1159), .A2(new_n839), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n1135), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1104), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1162), .A2(KEYINPUT122), .A3(new_n1165), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1089), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT109), .B1(G290), .B2(G1986), .ZN(new_n1171));
  NAND2_X1  g746(.A1(G290), .A2(G1986), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1171), .B(new_n1172), .Z(new_n1173));
  OAI21_X1  g748(.A(new_n978), .B1(new_n965), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n990), .B1(new_n1170), .B2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g750(.A1(new_n884), .A2(new_n886), .ZN(new_n1177));
  NOR4_X1   g751(.A1(G227), .A2(G229), .A3(new_n461), .A4(G401), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1177), .A2(new_n954), .A3(new_n1178), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


