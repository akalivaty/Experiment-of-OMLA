//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203,
    new_n1204, new_n1205, new_n1206;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  INV_X1    g0005(.A(KEYINPUT1), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G116), .A2(G270), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G87), .A2(G250), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G50), .B2(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n205), .B1(KEYINPUT65), .B2(new_n206), .C1(new_n216), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n205), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT64), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n222), .A2(new_n226), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n213), .A2(G1698), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G226), .B2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n251), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n225), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n250), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n248), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n218), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n268), .A2(new_n269), .ZN(new_n271));
  OAI21_X1  g0071(.A(G179), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G169), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n272), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n224), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT66), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(G77), .B1(G50), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n224), .B2(G68), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n225), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT11), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT12), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n224), .A3(G1), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n292), .B2(G68), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n294));
  INV_X1    g0094(.A(new_n286), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G1), .B2(new_n224), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n293), .B(new_n294), .C1(new_n217), .C2(new_n296), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT70), .Z(new_n298));
  NAND2_X1  g0098(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n288), .A2(KEYINPUT71), .A3(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n268), .B(new_n269), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(G190), .B1(new_n301), .B2(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n273), .A2(G200), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n278), .A2(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT8), .B(G58), .Z(new_n309));
  AOI22_X1  g0109(.A1(new_n281), .A2(new_n309), .B1(G150), .B2(new_n282), .ZN(new_n310));
  OAI21_X1  g0110(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G50), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n291), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n296), .A2(new_n313), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT9), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT3), .B(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G222), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G223), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n263), .C1(G77), .C2(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(new_n250), .ZN(new_n325));
  INV_X1    g0125(.A(G226), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n265), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n314), .A2(KEYINPUT9), .A3(new_n315), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n318), .A2(new_n328), .A3(new_n329), .A4(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT68), .B1(new_n332), .B2(KEYINPUT10), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(KEYINPUT10), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT68), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n332), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT10), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT67), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT67), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n332), .A2(new_n340), .A3(KEYINPUT10), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n333), .A2(new_n336), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n327), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n327), .A2(G179), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n316), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n309), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n279), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n349), .A2(new_n286), .B1(new_n350), .B2(new_n291), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n350), .B2(new_n296), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G232), .A2(G1698), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n321), .A2(G238), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n319), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n263), .C1(G107), .C2(new_n319), .ZN(new_n356));
  INV_X1    g0156(.A(G244), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n325), .C1(new_n357), .C2(new_n265), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(G179), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n343), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n352), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n308), .A2(new_n342), .A3(new_n346), .A4(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n256), .A2(G33), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT73), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n255), .A2(new_n257), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n368), .B2(new_n224), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT7), .B(new_n224), .C1(new_n363), .C2(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT74), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n258), .A2(new_n372), .A3(KEYINPUT7), .A4(new_n224), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n212), .A2(new_n217), .ZN(new_n376));
  OAI21_X1  g0176(.A(G20), .B1(new_n376), .B2(new_n201), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n282), .A2(G159), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(KEYINPUT16), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n319), .B2(G20), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n370), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n380), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n295), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n309), .A2(new_n291), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n296), .B2(new_n309), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n326), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n319), .B(new_n394), .C1(G223), .C2(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n262), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n325), .B1(new_n265), .B2(new_n213), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G169), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(G179), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT18), .B1(new_n393), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(G190), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n400), .A2(G200), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n389), .A2(new_n408), .A3(new_n392), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n410), .A2(new_n411), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n352), .B1(G200), .B2(new_n358), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n330), .B2(new_n358), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n407), .A2(new_n412), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n362), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G45), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G1), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT5), .B(G41), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n263), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G270), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n418), .A2(new_n249), .A3(G1), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n215), .A2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G257), .B2(G1698), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n262), .B1(new_n319), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G303), .B2(new_n319), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G179), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT21), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(G169), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G116), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n291), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n292), .B(new_n295), .C1(G1), .C2(new_n254), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G283), .ZN(new_n439));
  INV_X1    g0239(.A(G97), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n224), .C1(G33), .C2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n286), .C1(new_n224), .C2(G116), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT20), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n437), .B1(new_n436), .B2(new_n438), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n432), .A2(KEYINPUT79), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(G169), .A3(new_n429), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n435), .A2(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n429), .A2(G200), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n330), .C2(new_n429), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n319), .A2(new_n224), .A3(G87), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT22), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n254), .A2(G20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n224), .A2(G107), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT23), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT80), .B(KEYINPUT24), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n461), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n455), .A2(new_n457), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n286), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n438), .A2(new_n214), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n291), .A2(new_n214), .ZN(new_n468));
  XOR2_X1   g0268(.A(new_n468), .B(KEYINPUT25), .Z(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n319), .B1(G250), .B2(G1698), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n321), .A2(G257), .ZN(new_n472));
  INV_X1    g0272(.A(G294), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n471), .A2(new_n472), .B1(new_n254), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n263), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n421), .A2(G264), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n424), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G179), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n470), .B(new_n480), .C1(G169), .C2(new_n478), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n465), .A2(new_n467), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(G190), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(G200), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n482), .A2(new_n469), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n453), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n438), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G87), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n456), .A2(G97), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n224), .B1(new_n251), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n489), .A2(new_n490), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n319), .A2(new_n224), .A3(G68), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n286), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n348), .A2(new_n291), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n488), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n357), .A2(G1698), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n319), .B(new_n502), .C1(G238), .C2(G1698), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n262), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n262), .B(G250), .C1(G1), .C2(new_n418), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n505), .A2(new_n507), .A3(new_n423), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n500), .B(KEYINPUT77), .C1(new_n501), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT77), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n508), .A2(new_n501), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n488), .A2(new_n498), .A3(new_n499), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(G190), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n479), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n348), .B(KEYINPUT76), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n498), .B(new_n499), .C1(new_n438), .C2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(new_n518), .C1(G169), .C2(new_n508), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT78), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n515), .A2(KEYINPUT78), .A3(new_n519), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n292), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n440), .A2(new_n214), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(new_n492), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n384), .A2(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n295), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n525), .B(new_n533), .C1(G97), .C2(new_n487), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n319), .A2(G244), .A3(new_n321), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n319), .A2(KEYINPUT4), .A3(G244), .A4(new_n321), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n319), .A2(G250), .A3(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n537), .A2(new_n439), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n263), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n421), .A2(G257), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n424), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n543), .A2(new_n330), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n534), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n543), .A2(G179), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n533), .A2(new_n525), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n440), .B2(new_n438), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n343), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n417), .A2(new_n486), .A3(new_n524), .A4(new_n554), .ZN(G372));
  INV_X1    g0355(.A(new_n346), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n306), .A2(new_n307), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n305), .A2(G179), .B1(KEYINPUT72), .B2(KEYINPUT14), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n303), .B1(new_n558), .B2(new_n276), .ZN(new_n559));
  INV_X1    g0359(.A(new_n361), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n413), .A2(new_n412), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n407), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n563), .B2(new_n342), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n481), .A2(new_n449), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n546), .A2(new_n551), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n500), .B(new_n514), .C1(new_n501), .C2(new_n508), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n567), .A2(new_n485), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n551), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n522), .A2(KEYINPUT26), .A3(new_n523), .A4(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n519), .C1(new_n572), .C2(KEYINPUT81), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT26), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n519), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n551), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n572), .A2(KEYINPUT81), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n417), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n566), .A2(new_n578), .ZN(G369));
  AND2_X1   g0379(.A1(new_n485), .A2(new_n481), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n290), .A2(G20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n247), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n582), .A2(KEYINPUT27), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(KEYINPUT27), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(G213), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G343), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n449), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n587), .B(KEYINPUT84), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n481), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n446), .A2(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n453), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n449), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G330), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT83), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n470), .A2(new_n587), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n580), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n587), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n481), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n592), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT85), .ZN(G399));
  INV_X1    g0404(.A(new_n227), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(G41), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G1), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n492), .A2(new_n493), .A3(new_n436), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(new_n223), .B2(new_n607), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT28), .ZN(new_n611));
  INV_X1    g0411(.A(new_n590), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n573), .B2(new_n577), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT29), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n551), .A2(new_n575), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n619), .A2(KEYINPUT87), .A3(KEYINPUT26), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT87), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n522), .A2(new_n523), .A3(new_n571), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n574), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n570), .A2(new_n519), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n587), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT29), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n478), .A2(new_n542), .A3(new_n541), .ZN(new_n629));
  INV_X1    g0429(.A(new_n508), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n629), .A2(new_n431), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT30), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n430), .A2(G179), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n477), .A3(new_n630), .A4(new_n543), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n587), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT31), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n486), .A2(new_n554), .A3(new_n524), .A4(new_n612), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(KEYINPUT31), .A3(new_n590), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n618), .A2(new_n628), .B1(G330), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n611), .B1(new_n643), .B2(G1), .ZN(G364));
  NOR2_X1   g0444(.A1(new_n479), .A2(new_n501), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n224), .A2(new_n330), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G50), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n330), .A2(G179), .A3(G200), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n224), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n224), .A2(G190), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n479), .A3(new_n501), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT89), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G159), .ZN(new_n661));
  OAI221_X1 g0461(.A(new_n649), .B1(new_n440), .B2(new_n654), .C1(new_n661), .C2(KEYINPUT32), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT32), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n645), .A2(new_n655), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n258), .B1(new_n665), .B2(G68), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n501), .A2(G179), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n646), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G87), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n479), .A2(G200), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n646), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n655), .A2(new_n671), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n672), .A2(new_n212), .B1(new_n673), .B2(new_n350), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT88), .Z(new_n675));
  NAND4_X1  g0475(.A1(new_n663), .A2(new_n666), .A3(new_n670), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n655), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI211_X1 g0478(.A(new_n662), .B(new_n676), .C1(G107), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G311), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G322), .ZN(new_n682));
  OAI221_X1 g0482(.A(new_n258), .B1(new_n672), .B2(new_n682), .C1(new_n651), .C2(new_n473), .ZN(new_n683));
  AOI211_X1 g0483(.A(new_n681), .B(new_n683), .C1(G303), .C2(new_n669), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n660), .A2(G329), .ZN(new_n685));
  XNOR2_X1  g0485(.A(KEYINPUT33), .B(G317), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n665), .A2(new_n686), .B1(new_n678), .B2(G283), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(G326), .B2(new_n648), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT91), .Z(new_n691));
  AOI21_X1  g0491(.A(new_n225), .B1(G20), .B2(new_n343), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n608), .B1(G45), .B2(new_n581), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n319), .A2(G355), .A3(new_n227), .ZN(new_n695));
  INV_X1    g0495(.A(new_n368), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n605), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n418), .B2(new_n245), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n223), .A2(G45), .ZN(new_n699));
  OAI221_X1 g0499(.A(new_n695), .B1(G116), .B2(new_n227), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G13), .A2(G33), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G20), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n692), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n693), .A2(new_n694), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n596), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n703), .ZN(new_n708));
  INV_X1    g0508(.A(new_n598), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n694), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n706), .A2(new_n708), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(G396));
  NOR2_X1   g0513(.A1(new_n361), .A2(new_n587), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n352), .A2(new_n587), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n415), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n714), .B1(new_n716), .B2(new_n361), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n612), .B(new_n717), .C1(new_n573), .C2(new_n577), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n615), .A2(new_n617), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n642), .A2(G330), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n694), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n721), .A2(KEYINPUT93), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n692), .A2(new_n701), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n672), .ZN(new_n728));
  INV_X1    g0528(.A(new_n673), .ZN(new_n729));
  AOI22_X1  g0529(.A1(G143), .A2(new_n728), .B1(new_n729), .B2(G159), .ZN(new_n730));
  INV_X1    g0530(.A(G137), .ZN(new_n731));
  INV_X1    g0531(.A(G150), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n730), .B1(new_n731), .B2(new_n647), .C1(new_n732), .C2(new_n664), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n678), .A2(G68), .ZN(new_n735));
  INV_X1    g0535(.A(G132), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n696), .B(new_n735), .C1(new_n659), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(G50), .B2(new_n669), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n734), .B(new_n738), .C1(new_n212), .C2(new_n651), .ZN(new_n739));
  INV_X1    g0539(.A(new_n654), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n740), .A2(G97), .B1(G116), .B2(new_n729), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n665), .A2(G283), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n660), .A2(G311), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n258), .B1(new_n668), .B2(new_n214), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n647), .A2(new_n745), .B1(new_n677), .B2(new_n493), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n744), .B(new_n746), .C1(G294), .C2(new_n728), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n739), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n692), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n694), .B1(G77), .B2(new_n727), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT92), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n702), .B2(new_n717), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n725), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(G384));
  OAI211_X1 g0555(.A(new_n413), .B(new_n412), .C1(new_n404), .C2(new_n405), .ZN(new_n756));
  INV_X1    g0556(.A(new_n585), .ZN(new_n757));
  AOI21_X1  g0557(.A(G20), .B1(new_n365), .B2(new_n367), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n371), .B(new_n373), .C1(new_n758), .C2(KEYINPUT7), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n379), .B1(new_n759), .B2(G68), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT16), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n295), .B1(new_n760), .B2(KEYINPUT16), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n391), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n756), .A2(new_n757), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n401), .A2(new_n402), .A3(new_n585), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n379), .B1(new_n384), .B2(G68), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n286), .B1(new_n767), .B2(KEYINPUT16), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n760), .B2(KEYINPUT16), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n766), .B1(new_n769), .B2(new_n391), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT37), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n410), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT94), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n770), .A2(new_n410), .A3(KEYINPUT94), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT95), .ZN(new_n777));
  INV_X1    g0577(.A(new_n766), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n410), .B1(new_n763), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(KEYINPUT37), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n777), .B1(new_n776), .B2(new_n780), .ZN(new_n782));
  OAI211_X1 g0582(.A(KEYINPUT38), .B(new_n765), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n776), .A2(new_n780), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT97), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT38), .A4(new_n765), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n770), .A2(new_n410), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n776), .B1(new_n771), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n756), .A2(new_n393), .A3(new_n757), .ZN(new_n794));
  AOI21_X1  g0594(.A(KEYINPUT38), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n636), .A2(KEYINPUT31), .A3(new_n587), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n639), .A2(new_n640), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n278), .A2(new_n304), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n304), .A2(new_n587), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n800), .A2(new_n557), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n800), .B2(new_n601), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n799), .A2(new_n803), .A3(KEYINPUT40), .A4(new_n717), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n797), .A2(KEYINPUT100), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT100), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n795), .B1(new_n784), .B2(new_n790), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n804), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(KEYINPUT38), .B1(new_n788), .B2(new_n765), .ZN(new_n811));
  INV_X1    g0611(.A(new_n783), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT96), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n799), .A2(new_n803), .A3(new_n717), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n765), .B1(new_n781), .B2(new_n782), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT38), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT96), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n818), .A3(new_n783), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n813), .A2(new_n814), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT40), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n417), .A2(new_n799), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n810), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n710), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n810), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(G330), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n824), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n618), .A2(new_n628), .A3(new_n417), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n566), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n830), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n800), .A2(new_n587), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n817), .A2(KEYINPUT39), .A3(new_n783), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(new_n808), .C2(KEYINPUT39), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n308), .A2(new_n801), .B1(new_n559), .B2(new_n587), .ZN(new_n838));
  INV_X1    g0638(.A(new_n714), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n718), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n813), .A2(new_n840), .A3(new_n819), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n406), .A2(new_n585), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT98), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT98), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n836), .A2(new_n845), .A3(new_n842), .A4(new_n841), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n833), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n247), .B2(new_n581), .ZN(new_n850));
  OAI211_X1 g0650(.A(G20), .B(new_n260), .C1(new_n530), .C2(KEYINPUT35), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n436), .B(new_n851), .C1(KEYINPUT35), .C2(new_n530), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI21_X1  g0653(.A(G77), .B1(new_n212), .B2(new_n217), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n223), .A2(new_n854), .B1(G50), .B2(new_n217), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(G1), .A3(new_n290), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n850), .A2(new_n853), .A3(new_n856), .ZN(G367));
  AOI21_X1  g0657(.A(new_n247), .B1(new_n581), .B2(G45), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n589), .B(KEYINPUT104), .Z(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n602), .B2(new_n588), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT105), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n709), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n598), .A2(KEYINPUT105), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(new_n643), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n568), .B1(new_n534), .B2(new_n612), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n571), .A2(new_n590), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n592), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT44), .Z(new_n871));
  NOR2_X1   g0671(.A1(new_n592), .A2(new_n869), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT45), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n598), .A2(new_n602), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n871), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n876), .B(new_n877), .Z(new_n878));
  NAND2_X1  g0678(.A1(new_n866), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n643), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n606), .B(KEYINPUT41), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n859), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n869), .A2(new_n589), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  INV_X1    g0684(.A(new_n519), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n500), .A2(new_n601), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n575), .B2(new_n886), .ZN(new_n888));
  MUX2_X1   g0688(.A(new_n887), .B(new_n888), .S(KEYINPUT101), .Z(new_n889));
  XNOR2_X1  g0689(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n551), .B1(new_n867), .B2(new_n481), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n612), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n884), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT103), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n884), .A2(new_n893), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n891), .B1(KEYINPUT43), .B2(new_n889), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n874), .A2(new_n869), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n703), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n697), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n704), .B1(new_n227), .B2(new_n348), .C1(new_n904), .C2(new_n238), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n660), .A2(G317), .B1(G283), .B2(new_n729), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n906), .B1(new_n214), .B2(new_n651), .C1(new_n680), .C2(new_n647), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n368), .B1(new_n473), .B2(new_n664), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n672), .A2(new_n745), .B1(new_n677), .B2(new_n440), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n669), .A2(G116), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT46), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n740), .A2(G68), .B1(G143), .B2(new_n648), .ZN(new_n913));
  INV_X1    g0713(.A(G159), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(new_n664), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n319), .B1(new_n212), .B2(new_n668), .C1(new_n659), .C2(new_n731), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n313), .A2(new_n673), .B1(new_n677), .B2(new_n350), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n728), .A2(G150), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n910), .A2(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT47), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n694), .B(new_n905), .C1(new_n921), .C2(new_n750), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n882), .A2(new_n901), .B1(new_n903), .B2(new_n922), .ZN(G387));
  NAND2_X1  g0723(.A1(new_n865), .A2(new_n859), .ZN(new_n924));
  AOI22_X1  g0724(.A1(G322), .A2(new_n648), .B1(new_n665), .B2(G311), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n925), .B1(new_n745), .B2(new_n673), .C1(new_n926), .C2(new_n672), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT48), .ZN(new_n928));
  INV_X1    g0728(.A(G283), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n928), .B1(new_n929), .B2(new_n651), .C1(new_n473), .C2(new_n668), .ZN(new_n930));
  XNOR2_X1  g0730(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n660), .A2(G326), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n696), .B1(G116), .B2(new_n678), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n659), .A2(new_n732), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n665), .A2(new_n309), .ZN(new_n937));
  INV_X1    g0737(.A(new_n517), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n740), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n217), .B2(new_n673), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n669), .A2(G77), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n696), .B(new_n941), .C1(new_n914), .C2(new_n647), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n672), .A2(new_n313), .B1(new_n677), .B2(new_n440), .ZN(new_n943));
  OR4_X1    g0743(.A1(new_n937), .A2(new_n940), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n935), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n692), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n602), .A2(new_n902), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n697), .B1(new_n235), .B2(new_n418), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n319), .A2(new_n609), .A3(new_n227), .ZN(new_n949));
  AOI211_X1 g0749(.A(G45), .B(new_n609), .C1(G68), .C2(G77), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n309), .A2(new_n313), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT50), .Z(new_n952));
  AOI22_X1  g0752(.A1(new_n948), .A2(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n227), .A2(G107), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n704), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n946), .A2(new_n947), .A3(new_n694), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n606), .B1(new_n865), .B2(new_n643), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n924), .B(new_n956), .C1(new_n866), .C2(new_n957), .ZN(G393));
  NAND2_X1  g0758(.A1(new_n869), .A2(new_n703), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n704), .B1(new_n904), .B2(new_n242), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G97), .B2(new_n605), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n694), .B1(new_n961), .B2(KEYINPUT108), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n258), .B1(new_n677), .B2(new_n214), .C1(new_n929), .C2(new_n668), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n660), .B2(G322), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT109), .Z(new_n965));
  OAI22_X1  g0765(.A1(new_n647), .A2(new_n926), .B1(new_n672), .B2(new_n680), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT52), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n664), .A2(new_n745), .B1(new_n673), .B2(new_n473), .ZN(new_n968));
  INV_X1    g0768(.A(new_n651), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(G116), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT110), .Z(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n668), .A2(new_n217), .B1(new_n677), .B2(new_n493), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n696), .B1(new_n313), .B2(new_n664), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G143), .C2(new_n660), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n729), .A2(new_n309), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n740), .A2(G77), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n647), .A2(new_n732), .B1(new_n672), .B2(new_n914), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT51), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n750), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n962), .B(new_n981), .C1(KEYINPUT108), .C2(new_n961), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n878), .A2(new_n859), .B1(new_n959), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n866), .B(new_n878), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(new_n607), .ZN(G390));
  OAI21_X1  g0785(.A(new_n835), .B1(new_n808), .B2(KEYINPUT39), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n701), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n665), .A2(G107), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G116), .A2(new_n728), .B1(new_n729), .B2(G97), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n977), .A2(new_n258), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G294), .B2(new_n660), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n648), .A2(G283), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n991), .A2(new_n670), .A3(new_n735), .A4(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT114), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT54), .B(G143), .Z(new_n995));
  AOI22_X1  g0795(.A1(new_n665), .A2(G137), .B1(new_n729), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n740), .A2(G159), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT115), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G128), .A2(new_n648), .B1(new_n728), .B2(G132), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n669), .A2(G150), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT53), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n258), .B(new_n1002), .C1(G50), .C2(new_n678), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(G125), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n659), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n993), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n692), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n727), .A2(new_n309), .ZN(new_n1009));
  AND4_X1   g0809(.A1(new_n694), .A2(new_n987), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n716), .A2(new_n361), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n714), .B1(new_n627), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n838), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n834), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n840), .A2(new_n834), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1014), .A2(new_n797), .B1(new_n986), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n642), .A2(new_n803), .A3(G330), .A4(new_n717), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n799), .A2(G330), .A3(new_n717), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1018), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n803), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n1021), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(new_n1025), .B2(new_n1016), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1010), .B1(new_n1026), .B2(new_n859), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n566), .A2(new_n831), .A3(new_n828), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1019), .A2(new_n838), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT112), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1017), .A3(KEYINPUT112), .A4(new_n1012), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n717), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n838), .B1(new_n721), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1024), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n718), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n714), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1028), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1026), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1026), .A2(new_n1040), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n1042), .A3(new_n606), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1027), .B1(new_n1044), .B2(new_n1045), .ZN(G378));
  INV_X1    g0846(.A(KEYINPUT120), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1028), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n566), .A2(new_n831), .A3(KEYINPUT119), .A4(new_n828), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1026), .B2(new_n1040), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT118), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n316), .A2(new_n757), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n342), .A2(KEYINPUT116), .A3(new_n346), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT116), .B1(new_n342), .B2(new_n346), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n342), .A2(new_n346), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n1056), .A3(new_n1054), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1059), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1060), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n810), .A2(new_n825), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n810), .B2(new_n825), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n847), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1067), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n826), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n810), .A2(new_n825), .A3(new_n1067), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1072), .A2(new_n1073), .B1(new_n846), .B2(new_n844), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1053), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n846), .A3(new_n844), .A4(new_n1073), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1052), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1047), .B1(new_n1078), .B2(KEYINPUT57), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n847), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1052), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n607), .B1(new_n1081), .B2(KEYINPUT57), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1051), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1042), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT118), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1070), .A2(new_n1053), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT57), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(KEYINPUT120), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1079), .A2(new_n1082), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1067), .A2(new_n701), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n660), .A2(G283), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n696), .A2(G41), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n728), .A2(G107), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n941), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n740), .A2(G68), .B1(new_n938), .B2(new_n729), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n678), .A2(G58), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n440), .C2(new_n664), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1095), .B(new_n1098), .C1(G116), .C2(new_n648), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT58), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(G33), .A2(G41), .ZN(new_n1101));
  OR3_X1    g0901(.A1(new_n1093), .A2(G50), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n740), .A2(G150), .B1(G128), .B2(new_n728), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n647), .A2(new_n1005), .B1(new_n664), .B2(new_n736), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G137), .B2(new_n729), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n995), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1105), .C1(new_n668), .C2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT59), .ZN(new_n1108));
  INV_X1    g0908(.A(G124), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1101), .B1(new_n914), .B2(new_n677), .C1(new_n659), .C2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1102), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n692), .B1(new_n1100), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n726), .A2(new_n313), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1091), .A2(new_n694), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT117), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n859), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1090), .A2(new_n1117), .ZN(G375));
  INV_X1    g0918(.A(new_n1028), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1039), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n881), .ZN(new_n1122));
  OR3_X1    g0922(.A1(new_n1121), .A2(new_n1040), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n838), .A2(new_n701), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n694), .B1(G68), .B2(new_n727), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT121), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n440), .A2(new_n668), .B1(new_n664), .B2(new_n436), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n319), .B1(new_n678), .B2(G77), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n740), .A2(new_n938), .B1(KEYINPUT122), .B2(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(KEYINPUT122), .B2(new_n1128), .C1(new_n929), .C2(new_n672), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(G294), .C2(new_n648), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n214), .B2(new_n673), .C1(new_n745), .C2(new_n659), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT123), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n740), .A2(G50), .B1(G159), .B2(new_n669), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n736), .B2(new_n647), .C1(new_n664), .C2(new_n1106), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G137), .B2(new_n728), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n368), .B1(new_n660), .B2(G128), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n729), .A2(G150), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n1097), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1126), .B1(new_n1140), .B2(new_n692), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1120), .A2(new_n859), .B1(new_n1124), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1123), .A2(new_n1142), .ZN(G381));
  AND2_X1   g0943(.A1(new_n1043), .A2(new_n1027), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(G375), .A2(G384), .A3(G381), .A4(new_n1145), .ZN(new_n1146));
  OR2_X1    g0946(.A1(G387), .A2(G390), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1147), .A2(G396), .A3(G393), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(G407));
  NAND2_X1  g0949(.A1(new_n586), .A2(G213), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(G375), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(KEYINPUT124), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT124), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(G407), .A3(G213), .A4(new_n1153), .ZN(G409));
  NAND3_X1  g0954(.A1(new_n1090), .A2(G378), .A3(new_n1117), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n858), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1115), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1087), .B2(new_n1122), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1144), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1150), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n607), .B1(new_n1121), .B2(KEYINPUT60), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(KEYINPUT60), .C2(new_n1121), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1142), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n754), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT125), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(G384), .A3(new_n1142), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(G2897), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1150), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT125), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1171), .B1(new_n1174), .B2(new_n1169), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1161), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1173), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1160), .A2(new_n1150), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT62), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT61), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT62), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1160), .A2(new_n1182), .A3(new_n1150), .A4(new_n1178), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1177), .A2(new_n1180), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(G393), .B(G396), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(G387), .A2(G390), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT126), .B1(G387), .B2(G390), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1147), .A2(KEYINPUT126), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1160), .A2(KEYINPUT63), .A3(new_n1150), .A4(new_n1178), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1192), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n1181), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT63), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1175), .B1(new_n1160), .B2(new_n1150), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n1172), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1179), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1193), .A2(new_n1201), .ZN(G405));
  NAND2_X1  g1002(.A1(new_n1178), .A2(KEYINPUT127), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1192), .B(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1155), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G375), .B2(new_n1144), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1204), .B(new_n1206), .ZN(G402));
endmodule


