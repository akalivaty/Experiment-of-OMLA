//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT82), .ZN(new_n203));
  XNOR2_X1  g002(.A(G78gat), .B(G106gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT83), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n216), .A3(new_n211), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT76), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(new_n213), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n215), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n207), .B1(new_n225), .B2(KEYINPUT3), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n217), .A2(new_n213), .A3(new_n221), .A4(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n227), .A2(KEYINPUT78), .A3(new_n228), .A4(new_n215), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT29), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(KEYINPUT72), .ZN(new_n234));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236));
  INV_X1    g035(.A(G211gat), .ZN(new_n237));
  INV_X1    g036(.A(G218gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n234), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n228), .B1(new_n241), .B2(KEYINPUT29), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n227), .A2(KEYINPUT77), .A3(new_n215), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n242), .A2(new_n247), .A3(G228gat), .A4(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(G22gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(G228gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n241), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n230), .B2(new_n231), .ZN(new_n252));
  INV_X1    g051(.A(new_n225), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n240), .B2(new_n233), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n233), .B2(new_n240), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n255), .B2(new_n228), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n249), .B1(new_n248), .B2(new_n257), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n206), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT84), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n206), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n205), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n266), .A2(new_n258), .A3(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n260), .A2(new_n265), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n262), .A2(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n274), .A2(KEYINPUT66), .A3(new_n277), .A4(new_n275), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT24), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n280), .A2(new_n281), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n277), .A4(new_n275), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n289), .B1(new_n283), .B2(new_n285), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT28), .B1(new_n301), .B2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT26), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n273), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n275), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n302), .A2(new_n282), .A3(new_n305), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n299), .A2(KEYINPUT73), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n297), .B1(new_n292), .B2(new_n293), .ZN(new_n313));
  INV_X1    g112(.A(new_n310), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G226gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(KEYINPUT29), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n311), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n290), .A2(new_n288), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n321), .A2(new_n286), .B1(new_n278), .B2(new_n279), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT25), .B1(new_n322), .B2(new_n281), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT67), .B1(new_n323), .B2(new_n297), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n324), .A2(new_n326), .A3(new_n318), .A4(new_n310), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n241), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n315), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n318), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n310), .B1(new_n313), .B2(new_n325), .ZN(new_n332));
  AOI211_X1 g131(.A(KEYINPUT67), .B(new_n297), .C1(new_n292), .C2(new_n293), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n319), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n241), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT37), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337));
  INV_X1    g136(.A(new_n319), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n314), .B1(new_n299), .B2(KEYINPUT67), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n326), .ZN(new_n340));
  INV_X1    g139(.A(new_n318), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n311), .B2(new_n315), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n340), .A2(new_n342), .A3(new_n251), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n337), .B1(new_n343), .B2(new_n328), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT74), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n336), .B1(new_n346), .B2(KEYINPUT37), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G64gat), .ZN(new_n349));
  INV_X1    g148(.A(G92gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n272), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n353));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(G113gat), .ZN(new_n358));
  INV_X1    g157(.A(G120gat), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT1), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n362), .B(new_n360), .C1(new_n358), .C2(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n245), .A2(new_n366), .A3(new_n246), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n253), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT5), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n245), .A2(KEYINPUT3), .A3(new_n246), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n230), .A2(new_n374), .A3(new_n366), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT79), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n230), .A2(new_n374), .A3(new_n377), .A4(new_n366), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n372), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n368), .A2(new_n253), .A3(KEYINPUT80), .A4(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT4), .B1(new_n366), .B2(new_n225), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n366), .A2(new_n225), .A3(KEYINPUT4), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT80), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n380), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n373), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n383), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(new_n385), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n380), .A2(KEYINPUT5), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n391), .B(new_n393), .C1(new_n376), .C2(new_n378), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n357), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n391), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n396), .A3(new_n392), .ZN(new_n397));
  INV_X1    g196(.A(new_n357), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n372), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n376), .B2(new_n378), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n397), .B(new_n398), .C1(new_n401), .C2(new_n373), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n401), .B2(new_n373), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n329), .A2(new_n335), .A3(new_n351), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n351), .A2(new_n272), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n336), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n251), .B1(new_n340), .B2(new_n342), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT86), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n251), .C1(new_n340), .C2(new_n342), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n320), .A2(new_n327), .A3(new_n241), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n413), .A2(KEYINPUT37), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n410), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n270), .B1(new_n352), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n379), .A2(new_n396), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n380), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n371), .A2(new_n372), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(KEYINPUT39), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n398), .C1(KEYINPUT39), .C2(new_n422), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT40), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n425), .A2(new_n426), .B1(new_n357), .B2(new_n405), .ZN(new_n428));
  INV_X1    g227(.A(new_n407), .ZN(new_n429));
  INV_X1    g228(.A(new_n351), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n344), .A2(new_n430), .A3(new_n345), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n431), .B2(KEYINPUT30), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT30), .A4(new_n351), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT75), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n427), .B(new_n428), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n432), .A2(new_n434), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n404), .A2(new_n406), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n420), .A2(new_n435), .B1(new_n438), .B2(new_n270), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n366), .B1(new_n332), .B2(new_n333), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n324), .A2(new_n326), .A3(new_n368), .A4(new_n310), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(KEYINPUT71), .A3(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(G227gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(new_n317), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n447), .B(KEYINPUT64), .Z(new_n451));
  NOR3_X1   g250(.A1(new_n442), .A2(KEYINPUT34), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT70), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n442), .B2(new_n451), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  XOR2_X1   g257(.A(G71gat), .B(G99gat), .Z(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT69), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G15gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G43gat), .ZN(new_n462));
  INV_X1    g261(.A(G15gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n460), .B(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G43gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n458), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n455), .B1(new_n457), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n451), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n440), .B2(new_n441), .ZN(new_n471));
  NOR4_X1   g270(.A1(new_n471), .A2(new_n467), .A3(KEYINPUT70), .A4(new_n456), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n462), .A2(new_n466), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n471), .B2(KEYINPUT33), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT68), .B1(new_n471), .B2(new_n456), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n454), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n442), .A2(new_n451), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n457), .A2(new_n455), .A3(new_n468), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n475), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n476), .B1(new_n481), .B2(KEYINPUT32), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n471), .A2(KEYINPUT68), .A3(new_n456), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n452), .B1(new_n449), .B2(KEYINPUT34), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT36), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n480), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n480), .B2(new_n491), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n439), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n262), .A2(new_n264), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n268), .A2(new_n269), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n491), .A3(new_n480), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n500), .B2(new_n438), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n490), .B1(new_n485), .B2(new_n489), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n270), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  INV_X1    g304(.A(new_n437), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n506), .A2(new_n432), .A3(new_n434), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n496), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT11), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G169gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G197gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT12), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n515), .A2(new_n516), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT16), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n525), .A2(G1gat), .ZN(new_n530));
  OAI21_X1  g329(.A(G8gat), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n528), .B(new_n532), .C1(G1gat), .C2(new_n525), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n465), .A2(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(G50gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G43gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n537), .A3(KEYINPUT15), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n539), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n546), .B(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(new_n544), .A3(new_n542), .A4(new_n538), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT89), .B1(new_n536), .B2(G43gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n465), .A3(G50gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n554), .A3(new_n537), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT88), .B(KEYINPUT15), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n548), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n534), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT13), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n531), .A2(new_n533), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n558), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n534), .ZN(new_n568));
  OAI211_X1 g367(.A(KEYINPUT17), .B(new_n548), .C1(new_n551), .C2(new_n557), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n560), .B(new_n565), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n563), .B1(new_n573), .B2(KEYINPUT18), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n524), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n524), .A3(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(G71gat), .B2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n590), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n564), .B1(KEYINPUT21), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G183gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n534), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G183gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT93), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n597), .B2(new_n600), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n608), .A2(new_n610), .ZN(new_n613));
  OAI21_X1  g412(.A(G211gat), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n612), .A2(G211gat), .A3(new_n613), .ZN(new_n616));
  OAI22_X1  g415(.A1(new_n606), .A2(new_n607), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n600), .ZN(new_n618));
  INV_X1    g417(.A(new_n604), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n616), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n614), .A4(new_n605), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n632));
  AND2_X1   g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(G99gat), .A2(G106gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(KEYINPUT8), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT7), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G85gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n350), .ZN(new_n642));
  NAND3_X1  g441(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n637), .A2(new_n640), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n636), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n558), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n624), .A2(KEYINPUT41), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n637), .A2(new_n642), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n640), .A2(new_n643), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n636), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n635), .A3(new_n631), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n567), .A2(new_n569), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n567), .A2(KEYINPUT95), .A3(new_n569), .A4(new_n653), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AOI211_X1 g460(.A(new_n659), .B(new_n648), .C1(new_n656), .C2(new_n657), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n628), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n661), .ZN(new_n664));
  INV_X1    g463(.A(new_n662), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n627), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n623), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n644), .B1(new_n635), .B2(new_n631), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n586), .A2(new_n590), .A3(new_n588), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n590), .B1(new_n586), .B2(new_n588), .ZN(new_n671));
  OAI22_X1  g470(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n645), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n651), .A2(KEYINPUT96), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n674), .A3(new_n594), .ZN(new_n675));
  NAND2_X1  g474(.A1(G230gat), .A2(G233gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(G120gat), .B(G148gat), .Z(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT98), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT97), .B(G176gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n645), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n673), .A2(new_n675), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT10), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n678), .B(new_n683), .C1(new_n687), .C2(new_n677), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT99), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT10), .B1(new_n673), .B2(new_n675), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n676), .B1(new_n690), .B2(new_n684), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n678), .A4(new_n683), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n683), .B1(new_n691), .B2(new_n678), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT100), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n699), .B(new_n695), .C1(new_n689), .C2(new_n693), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AND4_X1   g502(.A1(new_n510), .A2(new_n580), .A3(new_n667), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n506), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G1gat), .ZN(G1324gat));
  INV_X1    g505(.A(new_n436), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT16), .B(G8gat), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n708), .A2(KEYINPUT42), .A3(new_n709), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n712), .B(new_n713), .C1(new_n532), .C2(new_n708), .ZN(G1325gat));
  NOR2_X1   g513(.A1(new_n502), .A2(new_n503), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n704), .A2(new_n463), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n493), .B2(new_n494), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT36), .B1(new_n502), .B2(new_n503), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n480), .A2(new_n491), .A3(new_n492), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(KEYINPUT101), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n704), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n716), .B1(new_n724), .B2(new_n463), .ZN(G1326gat));
  NAND2_X1  g524(.A1(new_n704), .A2(new_n270), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n722), .A2(new_n439), .B1(new_n501), .B2(new_n508), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n666), .A2(new_n663), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n510), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n702), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n573), .A2(KEYINPUT18), .ZN(new_n738));
  INV_X1    g537(.A(new_n563), .ZN(new_n739));
  AND4_X1   g538(.A1(new_n524), .A2(new_n738), .A3(new_n576), .A4(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n577), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n737), .A2(new_n741), .A3(new_n623), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n733), .A2(new_n506), .A3(new_n735), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n540), .B1(new_n743), .B2(KEYINPUT103), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT103), .B2(new_n743), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n741), .B1(new_n496), .B2(new_n509), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n732), .A2(new_n623), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n703), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n746), .A2(new_n540), .A3(new_n506), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n745), .A2(new_n751), .ZN(G1328gat));
  NAND4_X1  g551(.A1(new_n746), .A2(new_n541), .A3(new_n707), .A4(new_n749), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT46), .Z(new_n754));
  NAND2_X1  g553(.A1(new_n722), .A2(new_n439), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n509), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n731), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n757), .A2(new_n729), .B1(new_n510), .B2(new_n734), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n758), .A2(new_n707), .A3(new_n742), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n754), .B1(new_n541), .B2(new_n759), .ZN(G1329gat));
  INV_X1    g559(.A(new_n746), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n749), .A2(new_n465), .A3(new_n715), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n733), .A2(new_n723), .A3(new_n735), .A4(new_n742), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(G43gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n765), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n771), .ZN(G1330gat));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n536), .A3(new_n270), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n761), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n733), .A2(new_n270), .A3(new_n735), .A4(new_n742), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(G50gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n776), .A2(KEYINPUT105), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n776), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n778), .A2(new_n781), .ZN(G1331gat));
  INV_X1    g581(.A(new_n623), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n580), .A2(new_n731), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n737), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT106), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n785), .A2(KEYINPUT106), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n730), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n506), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n786), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n756), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n436), .B(new_n792), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1333gat));
  INV_X1    g594(.A(new_n715), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT108), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n788), .A2(new_n798), .A3(new_n715), .ZN(new_n799));
  INV_X1    g598(.A(G71gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n722), .A2(new_n800), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT107), .B1(new_n792), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n805), .A3(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT50), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n801), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1334gat));
  NAND2_X1  g611(.A1(new_n788), .A2(new_n270), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g613(.A1(new_n730), .A2(new_n732), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n741), .A2(new_n783), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT109), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT51), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NOR4_X1   g619(.A1(new_n730), .A2(new_n820), .A3(new_n732), .A4(new_n817), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n641), .A3(new_n506), .A4(new_n702), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n817), .A2(new_n703), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n758), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n506), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n826), .B2(new_n641), .ZN(G1336gat));
  INV_X1    g626(.A(new_n737), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(G92gat), .A3(new_n436), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n819), .B2(new_n821), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n733), .A2(new_n707), .A3(new_n735), .A4(new_n824), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G92gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n350), .B1(new_n831), .B2(KEYINPUT110), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n758), .A2(new_n836), .A3(new_n707), .A4(new_n824), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n834), .B1(new_n838), .B2(new_n840), .ZN(G1337gat));
  INV_X1    g640(.A(G99gat), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n822), .A2(new_n842), .A3(new_n715), .A4(new_n702), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n825), .A2(new_n723), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n842), .ZN(G1338gat));
  NOR3_X1   g644(.A1(new_n828), .A2(G106gat), .A3(new_n499), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT111), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n819), .B2(new_n821), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n733), .A2(new_n270), .A3(new_n735), .A4(new_n824), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G106gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1339gat));
  NAND4_X1  g654(.A1(new_n667), .A2(new_n698), .A3(new_n741), .A4(new_n701), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT112), .ZN(new_n857));
  INV_X1    g656(.A(new_n691), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n683), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n687), .A2(new_n677), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n691), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(KEYINPUT55), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n694), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n862), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n580), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(G229gat), .A3(G233gat), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n559), .A2(new_n562), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n871), .A2(new_n872), .B1(new_n518), .B2(new_n519), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n740), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n697), .B2(new_n700), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n731), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  AND4_X1   g675(.A1(new_n731), .A2(new_n865), .A3(new_n874), .A4(new_n868), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n783), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n500), .B1(new_n857), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n506), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(KEYINPUT114), .A3(new_n506), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n707), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n580), .A2(new_n358), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT115), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n880), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n436), .A3(new_n580), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT113), .B1(new_n889), .B2(G113gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(G1340gat));
  NAND2_X1  g691(.A1(new_n888), .A2(new_n436), .ZN(new_n893));
  OAI21_X1  g692(.A(G120gat), .B1(new_n893), .B2(new_n828), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT116), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n702), .A2(new_n359), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT117), .Z(new_n897));
  NAND2_X1  g696(.A1(new_n884), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1341gat));
  INV_X1    g698(.A(G127gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n900), .A3(new_n623), .ZN(new_n901));
  OAI21_X1  g700(.A(G127gat), .B1(new_n893), .B2(new_n783), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1342gat));
  NOR2_X1   g702(.A1(new_n732), .A2(G134gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n883), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT114), .B1(new_n879), .B2(new_n506), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n436), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n884), .A2(new_n909), .A3(new_n904), .ZN(new_n910));
  OAI21_X1  g709(.A(G134gat), .B1(new_n893), .B2(new_n732), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n908), .A2(new_n910), .A3(new_n914), .A4(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1343gat));
  AOI211_X1 g715(.A(new_n437), .B(new_n707), .C1(new_n718), .C2(new_n721), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n875), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n874), .B(KEYINPUT119), .C1(new_n697), .C2(new_n700), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT120), .B1(new_n866), .B2(new_n867), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n866), .A2(KEYINPUT120), .A3(new_n867), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n923), .A2(new_n580), .A3(new_n865), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n877), .B1(new_n926), .B2(new_n732), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT121), .B1(new_n927), .B2(new_n623), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n741), .A2(new_n864), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n931));
  AOI211_X1 g730(.A(new_n931), .B(KEYINPUT55), .C1(new_n860), .C2(new_n862), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n922), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n919), .A2(new_n875), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n731), .B1(new_n934), .B2(new_n921), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n929), .B(new_n783), .C1(new_n935), .C2(new_n877), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n928), .A2(new_n936), .A3(new_n857), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n270), .A2(KEYINPUT57), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n499), .B1(new_n857), .B2(new_n878), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n918), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n208), .B1(new_n945), .B2(new_n580), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n918), .A2(new_n942), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n208), .A3(new_n580), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT122), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT58), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n949), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT58), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n937), .A2(new_n939), .B1(new_n943), .B2(new_n942), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n953), .A2(new_n741), .A3(new_n918), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n951), .B(new_n952), .C1(new_n208), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n950), .A2(new_n955), .ZN(G1344gat));
  NAND3_X1  g755(.A1(new_n947), .A2(new_n209), .A3(new_n702), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n702), .B1(new_n917), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n960), .B1(new_n959), .B2(new_n917), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n857), .A2(new_n878), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n939), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n856), .B1(new_n927), .B2(new_n623), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT57), .B1(new_n964), .B2(new_n270), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n965), .B2(KEYINPUT124), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n967), .B(KEYINPUT57), .C1(new_n964), .C2(new_n270), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n961), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n958), .B1(new_n969), .B2(G148gat), .ZN(new_n970));
  AOI211_X1 g769(.A(KEYINPUT59), .B(new_n209), .C1(new_n945), .C2(new_n702), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n957), .B1(new_n970), .B2(new_n971), .ZN(G1345gat));
  AOI21_X1  g771(.A(G155gat), .B1(new_n947), .B2(new_n623), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n623), .A2(G155gat), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT125), .Z(new_n975));
  AOI21_X1  g774(.A(new_n973), .B1(new_n945), .B2(new_n975), .ZN(G1346gat));
  NAND3_X1  g775(.A1(new_n947), .A2(new_n220), .A3(new_n731), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n953), .A2(new_n732), .A3(new_n918), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n220), .ZN(G1347gat));
  NOR2_X1   g778(.A1(new_n436), .A2(new_n506), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n879), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n981), .A2(new_n741), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(new_n514), .ZN(G1348gat));
  OAI21_X1  g782(.A(G176gat), .B1(new_n981), .B2(new_n828), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n703), .A2(G176gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n981), .B2(new_n985), .ZN(G1349gat));
  NAND3_X1  g785(.A1(new_n879), .A2(new_n623), .A3(new_n980), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(new_n596), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n988), .B1(new_n300), .B2(new_n987), .ZN(new_n989));
  XOR2_X1   g788(.A(new_n989), .B(KEYINPUT60), .Z(G1350gat));
  NOR2_X1   g789(.A1(new_n981), .A2(new_n732), .ZN(new_n991));
  NAND2_X1  g790(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g792(.A(KEYINPUT61), .B(G190gat), .Z(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n991), .B2(new_n994), .ZN(G1351gat));
  AND2_X1   g794(.A1(new_n722), .A2(new_n980), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n941), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n580), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n966), .A2(new_n968), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n1000), .A2(new_n996), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n741), .A2(new_n516), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1352gat));
  NAND3_X1  g802(.A1(new_n1000), .A2(new_n737), .A3(new_n996), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G204gat), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n703), .A2(G204gat), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  OR3_X1    g806(.A1(new_n997), .A2(KEYINPUT126), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(KEYINPUT126), .B1(new_n997), .B2(new_n1007), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1008), .A2(KEYINPUT62), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(KEYINPUT62), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1005), .A2(new_n1012), .ZN(G1353gat));
  OAI211_X1 g812(.A(new_n623), .B(new_n996), .C1(new_n966), .C2(new_n968), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(G211gat), .ZN(new_n1015));
  XOR2_X1   g814(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n237), .A3(new_n623), .ZN(new_n1018));
  NOR2_X1   g817(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1014), .A2(G211gat), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(G1354gat));
  AOI21_X1  g820(.A(G218gat), .B1(new_n998), .B2(new_n731), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n732), .A2(new_n238), .ZN(new_n1023));
  AOI21_X1  g822(.A(new_n1022), .B1(new_n1001), .B2(new_n1023), .ZN(G1355gat));
endmodule


