

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803;

  INV_X1 U368 ( .A(n695), .ZN(n346) );
  INV_X1 U369 ( .A(n710), .ZN(n348) );
  AND2_X2 U370 ( .A1(n622), .A2(n621), .ZN(n655) );
  XNOR2_X1 U371 ( .A(n347), .B(n346), .ZN(G57) );
  NAND2_X1 U372 ( .A1(n357), .A2(n356), .ZN(n347) );
  XNOR2_X1 U373 ( .A(n349), .B(n348), .ZN(G60) );
  NAND2_X1 U374 ( .A1(n360), .A2(n359), .ZN(n349) );
  INV_X2 U375 ( .A(G953), .ZN(n796) );
  BUF_X1 U376 ( .A(G104), .Z(n428) );
  XOR2_X1 U377 ( .A(n704), .B(n703), .Z(n350) );
  AND2_X2 U378 ( .A1(n455), .A2(n441), .ZN(n437) );
  NOR2_X2 U379 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X2 U380 ( .A(n480), .B(KEYINPUT39), .ZN(n680) );
  XNOR2_X2 U381 ( .A(n659), .B(KEYINPUT42), .ZN(n801) );
  INV_X1 U382 ( .A(KEYINPUT80), .ZN(n370) );
  AND2_X1 U383 ( .A1(n367), .A2(n365), .ZN(n364) );
  AND2_X1 U384 ( .A1(n451), .A2(n449), .ZN(n672) );
  AND2_X1 U385 ( .A1(n475), .A2(n474), .ZN(n473) );
  NAND2_X1 U386 ( .A1(n743), .A2(n752), .ZN(n463) );
  NAND2_X1 U387 ( .A1(n370), .A2(KEYINPUT2), .ZN(n368) );
  AND2_X1 U388 ( .A1(n366), .A2(KEYINPUT80), .ZN(n365) );
  INV_X1 U389 ( .A(KEYINPUT77), .ZN(n394) );
  INV_X1 U390 ( .A(KEYINPUT46), .ZN(n392) );
  XOR2_X1 U391 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n580) );
  XNOR2_X1 U392 ( .A(G146), .B(G125), .ZN(n577) );
  INV_X1 U393 ( .A(KEYINPUT76), .ZN(n371) );
  INV_X1 U394 ( .A(KEYINPUT2), .ZN(n366) );
  INV_X1 U395 ( .A(KEYINPUT53), .ZN(n373) );
  XNOR2_X1 U396 ( .A(n374), .B(n373), .ZN(G75) );
  AND2_X1 U397 ( .A1(n353), .A2(n352), .ZN(n706) );
  AND2_X1 U398 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U399 ( .A(n376), .B(KEYINPUT113), .ZN(n375) );
  NAND2_X1 U400 ( .A1(n422), .A2(n421), .ZN(n376) );
  XNOR2_X1 U401 ( .A(n372), .B(n371), .ZN(n423) );
  NOR2_X1 U402 ( .A1(n364), .A2(n363), .ZN(n362) );
  OR2_X1 U403 ( .A1(KEYINPUT2), .A2(n795), .ZN(n736) );
  AND2_X1 U404 ( .A1(n795), .A2(n417), .ZN(n397) );
  NAND2_X1 U405 ( .A1(n369), .A2(n368), .ZN(n363) );
  XNOR2_X1 U406 ( .A(n627), .B(KEYINPUT45), .ZN(n652) );
  AND2_X1 U407 ( .A1(n385), .A2(n669), .ZN(n351) );
  AND2_X1 U408 ( .A1(n386), .A2(n668), .ZN(n385) );
  XNOR2_X1 U409 ( .A(n672), .B(n394), .ZN(n386) );
  OR2_X1 U410 ( .A1(n719), .A2(n450), .ZN(n449) );
  AND2_X1 U411 ( .A1(n602), .A2(n645), .ZN(n603) );
  XNOR2_X1 U412 ( .A(n377), .B(KEYINPUT71), .ZN(n654) );
  AND2_X1 U413 ( .A1(n473), .A2(n470), .ZN(n405) );
  XNOR2_X1 U414 ( .A(n465), .B(KEYINPUT38), .ZN(n753) );
  XNOR2_X1 U415 ( .A(n463), .B(n462), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n536), .B(n535), .ZN(n737) );
  XNOR2_X1 U417 ( .A(n743), .B(n597), .ZN(n645) );
  BUF_X1 U418 ( .A(n782), .Z(n354) );
  XNOR2_X1 U419 ( .A(n565), .B(n564), .ZN(n622) );
  XNOR2_X1 U420 ( .A(n557), .B(n544), .ZN(n476) );
  XNOR2_X1 U421 ( .A(n580), .B(n577), .ZN(n434) );
  XNOR2_X1 U422 ( .A(G122), .B(G107), .ZN(n496) );
  XNOR2_X1 U423 ( .A(KEYINPUT7), .B(G116), .ZN(n498) );
  XNOR2_X1 U424 ( .A(G113), .B(G143), .ZN(n559) );
  XNOR2_X1 U425 ( .A(G125), .B(G140), .ZN(n446) );
  NAND2_X1 U426 ( .A1(n395), .A2(n351), .ZN(n393) );
  INV_X1 U427 ( .A(n786), .ZN(n352) );
  XNOR2_X1 U428 ( .A(n705), .B(n350), .ZN(n353) );
  XNOR2_X2 U429 ( .A(n534), .B(n533), .ZN(n641) );
  XNOR2_X2 U430 ( .A(n666), .B(n665), .ZN(n719) );
  XNOR2_X1 U431 ( .A(n574), .B(n576), .ZN(n435) );
  XNOR2_X2 U432 ( .A(n491), .B(n490), .ZN(n574) );
  XNOR2_X2 U433 ( .A(n355), .B(n595), .ZN(n604) );
  NAND2_X1 U434 ( .A1(n412), .A2(n616), .ZN(n355) );
  INV_X1 U435 ( .A(n786), .ZN(n356) );
  XNOR2_X1 U436 ( .A(n694), .B(n358), .ZN(n357) );
  INV_X1 U437 ( .A(n693), .ZN(n358) );
  INV_X1 U438 ( .A(n786), .ZN(n359) );
  XNOR2_X1 U439 ( .A(n709), .B(n361), .ZN(n360) );
  INV_X1 U440 ( .A(n708), .ZN(n361) );
  NAND2_X1 U441 ( .A1(n736), .A2(n362), .ZN(n372) );
  INV_X1 U442 ( .A(n735), .ZN(n367) );
  NAND2_X1 U443 ( .A1(n735), .A2(n370), .ZN(n369) );
  NAND2_X1 U444 ( .A1(n375), .A2(n796), .ZN(n374) );
  XNOR2_X1 U445 ( .A(n403), .B(n484), .ZN(n638) );
  NAND2_X1 U446 ( .A1(n486), .A2(n485), .ZN(n403) );
  NAND2_X1 U447 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U448 ( .A(n737), .ZN(n380) );
  NAND2_X1 U449 ( .A1(n658), .A2(n382), .ZN(n381) );
  INV_X1 U450 ( .A(n644), .ZN(n382) );
  NAND2_X1 U451 ( .A1(n384), .A2(n383), .ZN(n390) );
  INV_X1 U452 ( .A(n803), .ZN(n383) );
  NOR2_X1 U453 ( .A1(n801), .A2(n392), .ZN(n384) );
  NAND2_X1 U454 ( .A1(n387), .A2(n392), .ZN(n391) );
  NAND2_X1 U455 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U456 ( .A(n801), .ZN(n388) );
  INV_X1 U457 ( .A(n803), .ZN(n389) );
  NAND2_X1 U458 ( .A1(n391), .A2(n390), .ZN(n395) );
  XNOR2_X2 U459 ( .A(n393), .B(n469), .ZN(n683) );
  NAND2_X1 U460 ( .A1(n398), .A2(n396), .ZN(n420) );
  NAND2_X1 U461 ( .A1(n400), .A2(n397), .ZN(n396) );
  NAND2_X1 U462 ( .A1(n399), .A2(n425), .ZN(n398) );
  NAND2_X1 U463 ( .A1(n400), .A2(n795), .ZN(n399) );
  XNOR2_X2 U464 ( .A(n689), .B(KEYINPUT83), .ZN(n795) );
  XNOR2_X2 U465 ( .A(n653), .B(KEYINPUT81), .ZN(n400) );
  NAND2_X2 U466 ( .A1(n604), .A2(n603), .ZN(n436) );
  XNOR2_X1 U467 ( .A(n634), .B(n429), .ZN(n704) );
  NAND2_X1 U468 ( .A1(n437), .A2(n459), .ZN(n439) );
  INV_X1 U469 ( .A(n738), .ZN(n401) );
  BUF_X1 U470 ( .A(n604), .Z(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n484), .ZN(n404) );
  NAND2_X1 U472 ( .A1(n473), .A2(n470), .ZN(n663) );
  BUF_X1 U473 ( .A(n652), .Z(n735) );
  XNOR2_X2 U474 ( .A(n419), .B(n691), .ZN(n779) );
  XNOR2_X1 U475 ( .A(KEYINPUT4), .B(G137), .ZN(n544) );
  NOR2_X1 U476 ( .A1(n645), .A2(n513), .ZN(n512) );
  XNOR2_X1 U477 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U478 ( .A(n493), .B(n492), .ZN(n573) );
  XNOR2_X1 U479 ( .A(G116), .B(G113), .ZN(n493) );
  XNOR2_X1 U480 ( .A(KEYINPUT3), .B(G119), .ZN(n492) );
  INV_X1 U481 ( .A(n686), .ZN(n427) );
  NOR2_X1 U482 ( .A1(G953), .A2(G237), .ZN(n556) );
  XOR2_X1 U483 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n560) );
  XNOR2_X1 U484 ( .A(n428), .B(G140), .ZN(n551) );
  NOR2_X1 U485 ( .A1(n506), .A2(KEYINPUT104), .ZN(n502) );
  NOR2_X1 U486 ( .A1(n643), .A2(n644), .ZN(n657) );
  NAND2_X1 U487 ( .A1(n458), .A2(n457), .ZN(n456) );
  OR2_X2 U488 ( .A1(n518), .A2(n515), .ZN(n743) );
  NAND2_X1 U489 ( .A1(n517), .A2(n457), .ZN(n516) );
  XNOR2_X1 U490 ( .A(n579), .B(n433), .ZN(n432) );
  INV_X1 U491 ( .A(KEYINPUT4), .ZN(n433) );
  NAND2_X1 U492 ( .A1(n654), .A2(n753), .ZN(n480) );
  INV_X1 U493 ( .A(KEYINPUT34), .ZN(n487) );
  NOR2_X1 U494 ( .A1(n673), .A2(n407), .ZN(n471) );
  XNOR2_X1 U495 ( .A(n435), .B(n573), .ZN(n634) );
  INV_X1 U496 ( .A(KEYINPUT47), .ZN(n450) );
  INV_X1 U497 ( .A(G237), .ZN(n549) );
  XNOR2_X1 U498 ( .A(KEYINPUT96), .B(KEYINPUT9), .ZN(n499) );
  AND2_X1 U499 ( .A1(n416), .A2(n426), .ZN(n425) );
  INV_X1 U500 ( .A(KEYINPUT48), .ZN(n469) );
  INV_X1 U501 ( .A(G472), .ZN(n517) );
  NAND2_X1 U502 ( .A1(G902), .A2(G472), .ZN(n519) );
  XNOR2_X1 U503 ( .A(n526), .B(n467), .ZN(n740) );
  XNOR2_X1 U504 ( .A(n468), .B(KEYINPUT92), .ZN(n467) );
  INV_X1 U505 ( .A(KEYINPUT21), .ZN(n468) );
  XNOR2_X1 U506 ( .A(n497), .B(n495), .ZN(n568) );
  XNOR2_X1 U507 ( .A(n496), .B(KEYINPUT97), .ZN(n495) );
  XNOR2_X1 U508 ( .A(n499), .B(n498), .ZN(n497) );
  NAND2_X1 U509 ( .A1(G234), .A2(G237), .ZN(n537) );
  INV_X1 U510 ( .A(KEYINPUT30), .ZN(n462) );
  NAND2_X1 U511 ( .A1(n673), .A2(n407), .ZN(n474) );
  XNOR2_X1 U512 ( .A(G101), .B(KEYINPUT5), .ZN(n545) );
  XNOR2_X1 U513 ( .A(n529), .B(n448), .ZN(n566) );
  INV_X1 U514 ( .A(KEYINPUT8), .ZN(n448) );
  XNOR2_X1 U515 ( .A(n411), .B(n481), .ZN(n444) );
  XNOR2_X1 U516 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n481) );
  XNOR2_X1 U517 ( .A(n482), .B(n530), .ZN(n443) );
  XNOR2_X1 U518 ( .A(G110), .B(G146), .ZN(n482) );
  XNOR2_X1 U519 ( .A(G119), .B(G128), .ZN(n530) );
  XNOR2_X1 U520 ( .A(n563), .B(n562), .ZN(n707) );
  XNOR2_X1 U521 ( .A(n561), .B(n406), .ZN(n562) );
  AND2_X1 U522 ( .A1(n796), .A2(G227), .ZN(n550) );
  XNOR2_X1 U523 ( .A(n454), .B(n453), .ZN(n452) );
  INV_X1 U524 ( .A(KEYINPUT28), .ZN(n453) );
  NAND2_X1 U525 ( .A1(n657), .A2(n743), .ZN(n454) );
  INV_X1 U526 ( .A(KEYINPUT0), .ZN(n489) );
  BUF_X1 U527 ( .A(n737), .Z(n466) );
  XNOR2_X1 U528 ( .A(n692), .B(KEYINPUT62), .ZN(n693) );
  XNOR2_X1 U529 ( .A(n445), .B(n442), .ZN(n782) );
  XNOR2_X1 U530 ( .A(n447), .B(n789), .ZN(n445) );
  XNOR2_X1 U531 ( .A(n444), .B(n443), .ZN(n442) );
  NAND2_X1 U532 ( .A1(n566), .A2(G221), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n707), .B(KEYINPUT59), .ZN(n708) );
  XNOR2_X1 U534 ( .A(n431), .B(n430), .ZN(n429) );
  XNOR2_X1 U535 ( .A(n434), .B(n432), .ZN(n431) );
  NOR2_X1 U536 ( .A1(n796), .A2(G952), .ZN(n786) );
  INV_X1 U537 ( .A(KEYINPUT40), .ZN(n478) );
  INV_X1 U538 ( .A(KEYINPUT35), .ZN(n484) );
  INV_X1 U539 ( .A(n610), .ZN(n485) );
  XOR2_X1 U540 ( .A(n560), .B(n559), .Z(n406) );
  XNOR2_X1 U541 ( .A(KEYINPUT72), .B(KEYINPUT19), .ZN(n407) );
  AND2_X1 U542 ( .A1(n440), .A2(n439), .ZN(n408) );
  XOR2_X1 U543 ( .A(n734), .B(KEYINPUT112), .Z(n409) );
  XOR2_X1 U544 ( .A(n670), .B(KEYINPUT78), .Z(n410) );
  XOR2_X1 U545 ( .A(G137), .B(KEYINPUT24), .Z(n411) );
  INV_X1 U546 ( .A(G902), .ZN(n457) );
  AND2_X1 U547 ( .A1(n594), .A2(n593), .ZN(n412) );
  AND2_X1 U548 ( .A1(n620), .A2(n658), .ZN(n413) );
  AND2_X1 U549 ( .A1(n408), .A2(n605), .ZN(n414) );
  NAND2_X1 U550 ( .A1(n690), .A2(n735), .ZN(n415) );
  INV_X1 U551 ( .A(KEYINPUT104), .ZN(n511) );
  INV_X1 U552 ( .A(KEYINPUT1), .ZN(n441) );
  NAND2_X1 U553 ( .A1(n686), .A2(n687), .ZN(n416) );
  AND2_X1 U554 ( .A1(n426), .A2(n687), .ZN(n417) );
  XNOR2_X2 U555 ( .A(n419), .B(n691), .ZN(n418) );
  NAND2_X2 U556 ( .A1(n420), .A2(n415), .ZN(n419) );
  NAND2_X1 U557 ( .A1(n440), .A2(n439), .ZN(n648) );
  NOR2_X1 U558 ( .A1(n769), .A2(n409), .ZN(n421) );
  NAND2_X1 U559 ( .A1(n423), .A2(n415), .ZN(n422) );
  XNOR2_X2 U560 ( .A(n424), .B(G134), .ZN(n569) );
  XNOR2_X1 U561 ( .A(n424), .B(n578), .ZN(n430) );
  XNOR2_X2 U562 ( .A(n543), .B(G128), .ZN(n424) );
  NAND2_X1 U563 ( .A1(n427), .A2(KEYINPUT65), .ZN(n426) );
  NAND2_X1 U564 ( .A1(n663), .A2(n591), .ZN(n477) );
  NAND2_X1 U565 ( .A1(n472), .A2(n471), .ZN(n470) );
  NAND2_X1 U566 ( .A1(n502), .A2(n509), .ZN(n500) );
  INV_X1 U567 ( .A(n510), .ZN(n506) );
  NAND2_X1 U568 ( .A1(n649), .A2(n738), .ZN(n494) );
  OR2_X2 U569 ( .A1(n770), .A2(n456), .ZN(n455) );
  NAND2_X1 U570 ( .A1(n640), .A2(n639), .ZN(n606) );
  NAND2_X1 U571 ( .A1(n402), .A2(n414), .ZN(n639) );
  XNOR2_X2 U572 ( .A(n436), .B(KEYINPUT32), .ZN(n640) );
  NAND2_X1 U573 ( .A1(n438), .A2(KEYINPUT1), .ZN(n440) );
  NAND2_X1 U574 ( .A1(n459), .A2(n455), .ZN(n438) );
  NAND2_X1 U575 ( .A1(n455), .A2(n459), .ZN(n658) );
  NAND2_X2 U576 ( .A1(n683), .A2(n523), .ZN(n689) );
  XNOR2_X2 U577 ( .A(n446), .B(KEYINPUT10), .ZN(n789) );
  INV_X1 U578 ( .A(n719), .ZN(n722) );
  NOR2_X1 U579 ( .A1(n671), .A2(n410), .ZN(n451) );
  NAND2_X1 U580 ( .A1(n452), .A2(n658), .ZN(n664) );
  INV_X1 U581 ( .A(n555), .ZN(n458) );
  AND2_X2 U582 ( .A1(n461), .A2(n460), .ZN(n459) );
  NAND2_X1 U583 ( .A1(n555), .A2(G902), .ZN(n460) );
  NAND2_X1 U584 ( .A1(n770), .A2(n555), .ZN(n461) );
  XNOR2_X2 U585 ( .A(n787), .B(n553), .ZN(n770) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n518) );
  NAND2_X1 U587 ( .A1(n464), .A2(n642), .ZN(n601) );
  INV_X1 U588 ( .A(n408), .ZN(n464) );
  NAND2_X1 U589 ( .A1(n638), .A2(n611), .ZN(n613) );
  XNOR2_X1 U590 ( .A(n488), .B(n487), .ZN(n486) );
  BUF_X2 U591 ( .A(n677), .Z(n465) );
  NOR2_X1 U592 ( .A1(n465), .A2(n673), .ZN(n510) );
  INV_X1 U593 ( .A(n677), .ZN(n472) );
  NAND2_X1 U594 ( .A1(n677), .A2(n407), .ZN(n475) );
  XNOR2_X2 U595 ( .A(n483), .B(KEYINPUT90), .ZN(n787) );
  XNOR2_X2 U596 ( .A(n569), .B(n476), .ZN(n483) );
  XNOR2_X2 U597 ( .A(n514), .B(G146), .ZN(n557) );
  XNOR2_X2 U598 ( .A(n477), .B(n489), .ZN(n616) );
  XNOR2_X2 U599 ( .A(n479), .B(n478), .ZN(n803) );
  NAND2_X1 U600 ( .A1(n680), .A2(n655), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n483), .B(n548), .ZN(n692) );
  NAND2_X1 U602 ( .A1(n732), .A2(n616), .ZN(n488) );
  NAND2_X1 U603 ( .A1(n616), .A2(n413), .ZN(n715) );
  XNOR2_X2 U604 ( .A(G110), .B(KEYINPUT88), .ZN(n490) );
  XNOR2_X2 U605 ( .A(G107), .B(G101), .ZN(n491) );
  XNOR2_X1 U606 ( .A(n494), .B(n650), .ZN(G27) );
  XNOR2_X1 U607 ( .A(n494), .B(KEYINPUT84), .ZN(n669) );
  AND2_X1 U608 ( .A1(n500), .A2(n501), .ZN(n505) );
  NAND2_X1 U609 ( .A1(n725), .A2(n502), .ZN(n501) );
  NAND2_X1 U610 ( .A1(n505), .A2(n503), .ZN(n647) );
  NAND2_X1 U611 ( .A1(n508), .A2(n504), .ZN(n503) );
  AND2_X1 U612 ( .A1(n512), .A2(n510), .ZN(n504) );
  NAND2_X1 U613 ( .A1(n507), .A2(n512), .ZN(n674) );
  INV_X1 U614 ( .A(n725), .ZN(n507) );
  NOR2_X1 U615 ( .A1(n725), .A2(n511), .ZN(n508) );
  INV_X1 U616 ( .A(n512), .ZN(n509) );
  INV_X1 U617 ( .A(n657), .ZN(n513) );
  XNOR2_X2 U618 ( .A(G131), .B(KEYINPUT68), .ZN(n514) );
  NAND2_X1 U619 ( .A1(n692), .A2(G472), .ZN(n520) );
  NOR2_X1 U620 ( .A1(n692), .A2(n516), .ZN(n515) );
  AND2_X1 U621 ( .A1(G214), .A2(n556), .ZN(n521) );
  XOR2_X1 U622 ( .A(n698), .B(n697), .Z(n522) );
  NOR2_X1 U623 ( .A1(n800), .A2(n682), .ZN(n523) );
  AND2_X1 U624 ( .A1(n625), .A2(n624), .ZN(n524) );
  INV_X1 U625 ( .A(KEYINPUT44), .ZN(n612) );
  INV_X1 U626 ( .A(KEYINPUT65), .ZN(n687) );
  XNOR2_X1 U627 ( .A(n354), .B(n781), .ZN(n783) );
  BUF_X1 U628 ( .A(n464), .Z(n738) );
  XNOR2_X1 U629 ( .A(n784), .B(n783), .ZN(n785) );
  XNOR2_X2 U630 ( .A(G902), .B(KEYINPUT15), .ZN(n684) );
  NAND2_X1 U631 ( .A1(G234), .A2(n684), .ZN(n525) );
  XNOR2_X1 U632 ( .A(KEYINPUT20), .B(n525), .ZN(n531) );
  NAND2_X1 U633 ( .A1(n531), .A2(G221), .ZN(n526) );
  INV_X1 U634 ( .A(KEYINPUT93), .ZN(n527) );
  XNOR2_X1 U635 ( .A(n740), .B(n527), .ZN(n593) );
  INV_X1 U636 ( .A(G953), .ZN(n528) );
  NAND2_X1 U637 ( .A1(G234), .A2(n528), .ZN(n529) );
  NOR2_X1 U638 ( .A1(n782), .A2(G902), .ZN(n534) );
  NAND2_X1 U639 ( .A1(n531), .A2(G217), .ZN(n532) );
  XNOR2_X1 U640 ( .A(n532), .B(KEYINPUT25), .ZN(n533) );
  NAND2_X1 U641 ( .A1(n593), .A2(n641), .ZN(n536) );
  INV_X1 U642 ( .A(KEYINPUT66), .ZN(n535) );
  XNOR2_X1 U643 ( .A(n537), .B(KEYINPUT14), .ZN(n538) );
  XNOR2_X1 U644 ( .A(KEYINPUT70), .B(n538), .ZN(n540) );
  NAND2_X1 U645 ( .A1(n540), .A2(G902), .ZN(n587) );
  OR2_X1 U646 ( .A1(n796), .A2(n587), .ZN(n539) );
  NOR2_X1 U647 ( .A1(G900), .A2(n539), .ZN(n542) );
  NAND2_X1 U648 ( .A1(G952), .A2(n540), .ZN(n768) );
  OR2_X1 U649 ( .A1(n768), .A2(G953), .ZN(n590) );
  INV_X1 U650 ( .A(n590), .ZN(n541) );
  NOR2_X1 U651 ( .A1(n542), .A2(n541), .ZN(n644) );
  XNOR2_X2 U652 ( .A(G143), .B(KEYINPUT74), .ZN(n543) );
  NAND2_X1 U653 ( .A1(n556), .A2(G210), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n573), .B(n547), .ZN(n548) );
  NAND2_X1 U656 ( .A1(n457), .A2(n549), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n581), .A2(G214), .ZN(n752) );
  XNOR2_X1 U658 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U659 ( .A(n574), .B(n552), .ZN(n553) );
  INV_X1 U660 ( .A(KEYINPUT69), .ZN(n554) );
  XNOR2_X1 U661 ( .A(n554), .B(G469), .ZN(n555) );
  XNOR2_X1 U662 ( .A(n557), .B(n521), .ZN(n558) );
  XNOR2_X1 U663 ( .A(n558), .B(n789), .ZN(n563) );
  XNOR2_X2 U664 ( .A(G122), .B(G104), .ZN(n575) );
  XNOR2_X1 U665 ( .A(n575), .B(KEYINPUT95), .ZN(n561) );
  NAND2_X1 U666 ( .A1(n707), .A2(n457), .ZN(n565) );
  XOR2_X1 U667 ( .A(KEYINPUT13), .B(G475), .Z(n564) );
  NAND2_X1 U668 ( .A1(G217), .A2(n566), .ZN(n567) );
  XNOR2_X1 U669 ( .A(n568), .B(n567), .ZN(n570) );
  XNOR2_X1 U670 ( .A(n569), .B(n570), .ZN(n698) );
  NAND2_X1 U671 ( .A1(n698), .A2(n457), .ZN(n572) );
  XOR2_X1 U672 ( .A(KEYINPUT98), .B(G478), .Z(n571) );
  XNOR2_X1 U673 ( .A(n572), .B(n571), .ZN(n621) );
  INV_X1 U674 ( .A(n621), .ZN(n592) );
  NAND2_X1 U675 ( .A1(n622), .A2(n592), .ZN(n610) );
  XNOR2_X1 U676 ( .A(n575), .B(KEYINPUT16), .ZN(n576) );
  XOR2_X1 U677 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n578) );
  NAND2_X1 U678 ( .A1(G224), .A2(n796), .ZN(n579) );
  NAND2_X1 U679 ( .A1(n704), .A2(n684), .ZN(n585) );
  NAND2_X1 U680 ( .A1(n581), .A2(G210), .ZN(n583) );
  INV_X1 U681 ( .A(KEYINPUT75), .ZN(n582) );
  XNOR2_X2 U682 ( .A(n585), .B(n584), .ZN(n677) );
  NOR2_X1 U683 ( .A1(n610), .A2(n465), .ZN(n586) );
  AND2_X1 U684 ( .A1(n654), .A2(n586), .ZN(n671) );
  XOR2_X1 U685 ( .A(n671), .B(G143), .Z(G45) );
  INV_X1 U686 ( .A(n752), .ZN(n673) );
  INV_X1 U687 ( .A(n587), .ZN(n588) );
  NOR2_X1 U688 ( .A1(n796), .A2(G898), .ZN(n635) );
  NAND2_X1 U689 ( .A1(n588), .A2(n635), .ZN(n589) );
  NAND2_X1 U690 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U691 ( .A1(n622), .A2(n592), .ZN(n755) );
  INV_X1 U692 ( .A(n755), .ZN(n594) );
  INV_X1 U693 ( .A(KEYINPUT22), .ZN(n595) );
  INV_X1 U694 ( .A(KEYINPUT99), .ZN(n596) );
  XNOR2_X1 U695 ( .A(n596), .B(KEYINPUT6), .ZN(n597) );
  AND2_X1 U696 ( .A1(n402), .A2(n645), .ZN(n599) );
  AND2_X1 U697 ( .A1(n401), .A2(n641), .ZN(n598) );
  NAND2_X1 U698 ( .A1(n599), .A2(n598), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(G101), .ZN(G3) );
  INV_X1 U700 ( .A(KEYINPUT100), .ZN(n600) );
  XNOR2_X1 U701 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X1 U702 ( .A1(n743), .A2(n641), .ZN(n605) );
  XNOR2_X1 U703 ( .A(n606), .B(KEYINPUT85), .ZN(n611) );
  NAND2_X1 U704 ( .A1(n648), .A2(n737), .ZN(n614) );
  XNOR2_X1 U705 ( .A(n614), .B(KEYINPUT101), .ZN(n608) );
  INV_X1 U706 ( .A(n645), .ZN(n607) );
  NAND2_X1 U707 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U708 ( .A(n609), .B(KEYINPUT33), .ZN(n732) );
  XNOR2_X1 U709 ( .A(n613), .B(n612), .ZN(n626) );
  INV_X1 U710 ( .A(n614), .ZN(n615) );
  AND2_X1 U711 ( .A1(n615), .A2(n743), .ZN(n747) );
  NAND2_X1 U712 ( .A1(n616), .A2(n747), .ZN(n618) );
  XOR2_X1 U713 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n617) );
  XNOR2_X1 U714 ( .A(n618), .B(n617), .ZN(n729) );
  INV_X1 U715 ( .A(n743), .ZN(n619) );
  AND2_X1 U716 ( .A1(n466), .A2(n619), .ZN(n620) );
  NAND2_X1 U717 ( .A1(n729), .A2(n715), .ZN(n623) );
  NOR2_X1 U718 ( .A1(n622), .A2(n621), .ZN(n718) );
  NOR2_X1 U719 ( .A1(n655), .A2(n718), .ZN(n757) );
  XNOR2_X1 U720 ( .A(n757), .B(KEYINPUT79), .ZN(n660) );
  NAND2_X1 U721 ( .A1(n623), .A2(n660), .ZN(n625) );
  NAND2_X1 U722 ( .A1(n626), .A2(n524), .ZN(n627) );
  NAND2_X1 U723 ( .A1(n735), .A2(n796), .ZN(n633) );
  XOR2_X1 U724 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n629) );
  NAND2_X1 U725 ( .A1(G224), .A2(G953), .ZN(n628) );
  XNOR2_X1 U726 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U727 ( .A(KEYINPUT123), .B(n630), .ZN(n631) );
  NAND2_X1 U728 ( .A1(n631), .A2(G898), .ZN(n632) );
  NAND2_X1 U729 ( .A1(n633), .A2(n632), .ZN(n637) );
  NOR2_X1 U730 ( .A1(n634), .A2(n635), .ZN(n636) );
  XNOR2_X1 U731 ( .A(n637), .B(n636), .ZN(G69) );
  XNOR2_X1 U732 ( .A(n404), .B(G122), .ZN(G24) );
  XNOR2_X1 U733 ( .A(n639), .B(G110), .ZN(G12) );
  XNOR2_X1 U734 ( .A(n640), .B(G119), .ZN(G21) );
  INV_X1 U735 ( .A(n641), .ZN(n642) );
  NAND2_X1 U736 ( .A1(n740), .A2(n642), .ZN(n643) );
  XOR2_X2 U737 ( .A(KEYINPUT102), .B(n655), .Z(n725) );
  XOR2_X1 U738 ( .A(KEYINPUT105), .B(KEYINPUT36), .Z(n646) );
  XNOR2_X1 U739 ( .A(n647), .B(n646), .ZN(n649) );
  XOR2_X1 U740 ( .A(G125), .B(KEYINPUT37), .Z(n650) );
  INV_X1 U741 ( .A(n684), .ZN(n651) );
  NAND2_X1 U742 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U743 ( .A1(n753), .A2(n752), .ZN(n756) );
  NOR2_X1 U744 ( .A1(n755), .A2(n756), .ZN(n656) );
  XNOR2_X1 U745 ( .A(KEYINPUT41), .B(n656), .ZN(n751) );
  NOR2_X1 U746 ( .A1(n751), .A2(n664), .ZN(n659) );
  INV_X1 U747 ( .A(n660), .ZN(n662) );
  XOR2_X1 U748 ( .A(KEYINPUT67), .B(KEYINPUT47), .Z(n661) );
  NOR2_X1 U749 ( .A1(n662), .A2(n661), .ZN(n667) );
  NOR2_X2 U750 ( .A1(n664), .A2(n405), .ZN(n666) );
  INV_X1 U751 ( .A(KEYINPUT73), .ZN(n665) );
  NAND2_X1 U752 ( .A1(n667), .A2(n719), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n757), .A2(KEYINPUT47), .ZN(n670) );
  NOR2_X1 U754 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n675), .A2(n401), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n676), .B(KEYINPUT43), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n678), .A2(n465), .ZN(n679) );
  XNOR2_X1 U758 ( .A(n679), .B(KEYINPUT103), .ZN(n800) );
  BUF_X1 U759 ( .A(n680), .Z(n681) );
  NAND2_X1 U760 ( .A1(n681), .A2(n718), .ZN(n731) );
  INV_X1 U761 ( .A(n731), .ZN(n682) );
  XOR2_X1 U762 ( .A(KEYINPUT82), .B(n684), .Z(n685) );
  NAND2_X1 U763 ( .A1(n685), .A2(KEYINPUT2), .ZN(n686) );
  INV_X1 U764 ( .A(KEYINPUT2), .ZN(n688) );
  NOR2_X1 U765 ( .A1(n689), .A2(n688), .ZN(n690) );
  INV_X1 U766 ( .A(KEYINPUT64), .ZN(n691) );
  NAND2_X1 U767 ( .A1(n779), .A2(G472), .ZN(n694) );
  XOR2_X1 U768 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n695) );
  NAND2_X1 U769 ( .A1(n418), .A2(G478), .ZN(n699) );
  XNOR2_X1 U770 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n697) );
  XNOR2_X1 U771 ( .A(n699), .B(n522), .ZN(n701) );
  INV_X1 U772 ( .A(n786), .ZN(n700) );
  XNOR2_X1 U773 ( .A(n702), .B(KEYINPUT120), .ZN(G63) );
  NAND2_X1 U774 ( .A1(n418), .A2(G210), .ZN(n705) );
  XNOR2_X1 U775 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n703) );
  XNOR2_X1 U776 ( .A(n706), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U777 ( .A1(n779), .A2(G475), .ZN(n709) );
  XOR2_X1 U778 ( .A(KEYINPUT117), .B(KEYINPUT60), .Z(n710) );
  NOR2_X1 U779 ( .A1(n725), .A2(n715), .ZN(n712) );
  XOR2_X1 U780 ( .A(n428), .B(n712), .Z(G6) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n714) );
  XNOR2_X1 U782 ( .A(G107), .B(KEYINPUT106), .ZN(n713) );
  XNOR2_X1 U783 ( .A(n714), .B(n713), .ZN(n717) );
  INV_X1 U784 ( .A(n718), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n728), .A2(n715), .ZN(n716) );
  XOR2_X1 U786 ( .A(n717), .B(n716), .Z(G9) );
  XOR2_X1 U787 ( .A(G128), .B(KEYINPUT29), .Z(n721) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U789 ( .A(n721), .B(n720), .ZN(G30) );
  NOR2_X1 U790 ( .A1(n725), .A2(n722), .ZN(n724) );
  XNOR2_X1 U791 ( .A(G146), .B(KEYINPUT107), .ZN(n723) );
  XNOR2_X1 U792 ( .A(n724), .B(n723), .ZN(G48) );
  NOR2_X1 U793 ( .A1(n725), .A2(n729), .ZN(n726) );
  XOR2_X1 U794 ( .A(KEYINPUT108), .B(n726), .Z(n727) );
  XNOR2_X1 U795 ( .A(G113), .B(n727), .ZN(G15) );
  NOR2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U797 ( .A(G116), .B(n730), .Z(G18) );
  XNOR2_X1 U798 ( .A(G134), .B(n731), .ZN(G36) );
  INV_X1 U799 ( .A(n751), .ZN(n733) );
  BUF_X1 U800 ( .A(n732), .Z(n761) );
  NAND2_X1 U801 ( .A1(n733), .A2(n761), .ZN(n734) );
  NOR2_X1 U802 ( .A1(n738), .A2(n466), .ZN(n739) );
  XNOR2_X1 U803 ( .A(n739), .B(KEYINPUT50), .ZN(n746) );
  NOR2_X1 U804 ( .A1(n740), .A2(n641), .ZN(n741) );
  XOR2_X1 U805 ( .A(KEYINPUT49), .B(n741), .Z(n742) );
  NOR2_X1 U806 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U807 ( .A(KEYINPUT109), .B(n744), .ZN(n745) );
  NOR2_X1 U808 ( .A1(n746), .A2(n745), .ZN(n748) );
  NOR2_X1 U809 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U810 ( .A(KEYINPUT51), .B(n749), .Z(n750) );
  NOR2_X1 U811 ( .A1(n751), .A2(n750), .ZN(n764) );
  NOR2_X1 U812 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U813 ( .A1(n755), .A2(n754), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U815 ( .A(n758), .B(KEYINPUT110), .ZN(n759) );
  OR2_X1 U816 ( .A1(n760), .A2(n759), .ZN(n762) );
  AND2_X1 U817 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U818 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U819 ( .A(n765), .B(KEYINPUT111), .Z(n766) );
  XNOR2_X1 U820 ( .A(KEYINPUT52), .B(n766), .ZN(n767) );
  NOR2_X1 U821 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U822 ( .A1(n780), .A2(G469), .ZN(n777) );
  BUF_X1 U823 ( .A(n770), .Z(n775) );
  XNOR2_X1 U824 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n771) );
  XNOR2_X1 U825 ( .A(n771), .B(KEYINPUT114), .ZN(n772) );
  XOR2_X1 U826 ( .A(n772), .B(KEYINPUT58), .Z(n773) );
  XOR2_X1 U827 ( .A(n773), .B(KEYINPUT57), .Z(n774) );
  XNOR2_X1 U828 ( .A(n775), .B(n774), .ZN(n776) );
  XNOR2_X1 U829 ( .A(n777), .B(n776), .ZN(n778) );
  NOR2_X1 U830 ( .A1(n786), .A2(n778), .ZN(G54) );
  BUF_X1 U831 ( .A(n779), .Z(n780) );
  NAND2_X1 U832 ( .A1(n780), .A2(G217), .ZN(n784) );
  XOR2_X1 U833 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n781) );
  NOR2_X1 U834 ( .A1(n786), .A2(n785), .ZN(G66) );
  BUF_X1 U835 ( .A(n787), .Z(n788) );
  XNOR2_X1 U836 ( .A(n789), .B(n788), .ZN(n794) );
  XOR2_X1 U837 ( .A(G227), .B(n794), .Z(n790) );
  NAND2_X1 U838 ( .A1(n790), .A2(G900), .ZN(n791) );
  XOR2_X1 U839 ( .A(KEYINPUT125), .B(n791), .Z(n792) );
  NAND2_X1 U840 ( .A1(G953), .A2(n792), .ZN(n793) );
  XNOR2_X1 U841 ( .A(n793), .B(KEYINPUT126), .ZN(n799) );
  XNOR2_X1 U842 ( .A(n795), .B(n794), .ZN(n797) );
  NAND2_X1 U843 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U844 ( .A1(n799), .A2(n798), .ZN(G72) );
  XOR2_X1 U845 ( .A(G140), .B(n800), .Z(G42) );
  XNOR2_X1 U846 ( .A(G137), .B(KEYINPUT127), .ZN(n802) );
  XNOR2_X1 U847 ( .A(n802), .B(n801), .ZN(G39) );
  XOR2_X1 U848 ( .A(n803), .B(G131), .Z(G33) );
endmodule

