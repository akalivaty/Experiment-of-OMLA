//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n637,
    new_n640, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G235), .A2(G236), .A3(G237), .A4(G238), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT71), .B1(new_n469), .B2(G101), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  AOI211_X1 g047(.A(new_n471), .B(new_n472), .C1(new_n467), .C2(new_n468), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n464), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  INV_X1    g054(.A(new_n462), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n489), .B2(new_n490), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n501), .C1(new_n490), .C2(new_n489), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT5), .A4(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(KEYINPUT73), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(KEYINPUT74), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n512), .A2(new_n515), .A3(G62), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n504), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(G543), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(G543), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n526));
  INV_X1    g101(.A(new_n507), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT75), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n533), .B1(new_n530), .B2(new_n522), .C1(new_n528), .C2(new_n529), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT7), .Z(new_n536));
  XOR2_X1   g111(.A(KEYINPUT6), .B(G651), .Z(new_n537));
  OAI21_X1  g112(.A(G543), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n537), .B1(new_n540), .B2(new_n507), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n536), .B1(new_n541), .B2(G89), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n532), .A2(new_n534), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  INV_X1    g119(.A(new_n522), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT76), .B(G52), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OAI221_X1 g124(.A(new_n547), .B1(new_n519), .B2(new_n548), .C1(new_n549), .C2(new_n504), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n512), .A2(G56), .ZN(new_n553));
  AND2_X1   g128(.A1(G68), .A2(G543), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n552), .B(G651), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n554), .B1(new_n512), .B2(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT77), .B1(new_n556), .B2(new_n504), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n541), .A2(G81), .B1(new_n545), .B2(G43), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n528), .C2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n568), .B1(new_n540), .B2(new_n507), .ZN(new_n570));
  INV_X1    g145(.A(new_n567), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n572), .A3(G651), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n522), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n518), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n576), .A2(new_n578), .B1(new_n541), .B2(G91), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n574), .B1(new_n573), .B2(new_n579), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G166), .ZN(G303));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT80), .B1(new_n519), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n541), .A2(new_n587), .A3(G87), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n586), .A2(new_n588), .B1(G49), .B2(new_n545), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n540), .A2(new_n591), .A3(new_n507), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n590), .B1(new_n592), .B2(G651), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n590), .A3(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n589), .A2(new_n596), .ZN(G288));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT83), .B1(new_n519), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n541), .A2(new_n600), .A3(G86), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n512), .A2(G61), .ZN(new_n604));
  AND2_X1   g179(.A1(G73), .A2(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(G651), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n545), .A2(G48), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n605), .B1(new_n512), .B2(G61), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT82), .B1(new_n608), .B2(new_n504), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n602), .A2(new_n606), .A3(new_n607), .A4(new_n609), .ZN(G305));
  AND2_X1   g185(.A1(new_n512), .A2(G60), .ZN(new_n611));
  AND2_X1   g186(.A1(G72), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT84), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(KEYINPUT84), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n541), .A2(G85), .B1(new_n545), .B2(G47), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT87), .B(G66), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n512), .A2(new_n619), .B1(G79), .B2(G543), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(new_n504), .ZN(new_n621));
  INV_X1    g196(.A(G54), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n522), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n522), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n519), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n541), .A2(G92), .A3(new_n626), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n621), .A2(new_n625), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n618), .B1(new_n632), .B2(G868), .ZN(G284));
  OAI21_X1  g208(.A(new_n618), .B1(new_n632), .B2(G868), .ZN(G321));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NOR2_X1   g210(.A1(G286), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G299), .B(KEYINPUT88), .Z(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n635), .ZN(G297));
  AOI21_X1  g213(.A(new_n636), .B1(new_n637), .B2(new_n635), .ZN(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n632), .B1(new_n640), .B2(G860), .ZN(G148));
  NOR2_X1   g216(.A1(new_n560), .A2(G868), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n632), .A2(new_n640), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(G868), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT89), .Z(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n469), .A2(new_n462), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT13), .Z(new_n649));
  INV_X1    g224(.A(G2100), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n481), .A2(G135), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n483), .A2(G123), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n463), .A2(G111), .ZN(new_n655));
  OAI21_X1  g230(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n651), .A2(new_n652), .A3(new_n659), .ZN(G156));
  XOR2_X1   g235(.A(G2427), .B(G2430), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT92), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT91), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT90), .B(KEYINPUT14), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(KEYINPUT93), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(KEYINPUT93), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  OAI22_X1  g244(.A1(new_n668), .A2(new_n669), .B1(new_n662), .B2(new_n665), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2451), .B(G2454), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G14), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n676), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G401));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT17), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(new_n650), .ZN(new_n688));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n684), .B2(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(new_n658), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(new_n703), .B(new_n702), .S(new_n695), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(G229));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n483), .B2(G129), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n469), .A2(G105), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n481), .A2(G141), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(G32), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n725));
  NAND2_X1  g300(.A1(G286), .A2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G21), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n719), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  AOI22_X1  g308(.A1(G128), .A2(new_n483), .B1(new_n481), .B2(G140), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(G116), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT99), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2067), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR4_X1   g317(.A1(new_n724), .A2(new_n725), .A3(new_n731), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n632), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G4), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1348), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n729), .A2(new_n730), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  NOR2_X1   g326(.A1(new_n657), .A2(new_n719), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT30), .B(G28), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n751), .B(new_n752), .C1(new_n719), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G27), .A2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G164), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n758), .C1(new_n721), .C2(new_n722), .ZN(new_n759));
  AND2_X1   g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n719), .B1(KEYINPUT24), .B2(G34), .ZN(new_n761));
  OAI22_X1  g336(.A1(G160), .A2(new_n719), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n759), .B1(G2084), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n727), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n727), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n719), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n719), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n766), .B1(new_n769), .B2(G2090), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n743), .A2(new_n750), .A3(new_n763), .A4(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT100), .B(KEYINPUT25), .Z(new_n772));
  NAND3_X1  g347(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n481), .A2(G139), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n774), .B(new_n775), .C1(new_n463), .C2(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G33), .B(new_n777), .S(G29), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT101), .ZN(new_n779));
  INV_X1    g354(.A(G2072), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT102), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n560), .A2(new_n727), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n727), .B2(G19), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n782), .B1(G1341), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G299), .A2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n727), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n769), .A2(G2090), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G1961), .B2(new_n765), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n785), .A2(G1341), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n762), .A2(G2084), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n779), .B2(new_n780), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n771), .A2(new_n786), .A3(new_n791), .A4(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G6), .B(G305), .S(G16), .Z(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT32), .B(G1981), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n545), .A2(G49), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n587), .B1(new_n541), .B2(G87), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n587), .A2(new_n512), .A3(G87), .A4(new_n518), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n595), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n593), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n589), .A2(KEYINPUT98), .A3(new_n596), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT33), .B(G1976), .Z(new_n817));
  OR2_X1    g392(.A1(G16), .A2(G23), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n817), .B1(new_n816), .B2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n727), .A2(G22), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n727), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1971), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT34), .B1(new_n805), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT34), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n804), .A2(new_n828), .A3(new_n824), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n719), .A2(G25), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n481), .A2(G131), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n483), .A2(G119), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n463), .A2(G107), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT94), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n830), .B1(new_n837), .B2(new_n719), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G1991), .Z(new_n839));
  XOR2_X1   g414(.A(new_n838), .B(new_n839), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n727), .A2(G24), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT95), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G290), .B2(G16), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(G1986), .Z(new_n844));
  NOR2_X1   g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n829), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT36), .B1(new_n827), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n826), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n799), .B1(new_n847), .B2(new_n850), .ZN(G311));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n798), .ZN(G150));
  NAND2_X1  g428(.A1(new_n632), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n504), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n519), .A2(new_n858), .B1(new_n859), .B2(new_n522), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n559), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n861), .A2(new_n555), .A3(new_n557), .A4(new_n558), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n855), .B(new_n865), .Z(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n861), .A2(new_n868), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  NAND2_X1  g448(.A1(new_n483), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n463), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G142), .B2(new_n481), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n648), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n777), .A2(KEYINPUT104), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n718), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n739), .B(G164), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n836), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n478), .B(new_n657), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n487), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n884), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n885), .B2(new_n888), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(G395));
  XNOR2_X1  g470(.A(G290), .B(G305), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n815), .A2(G303), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n813), .A2(new_n814), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(G166), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT107), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(KEYINPUT108), .Z(new_n909));
  OAI21_X1  g484(.A(new_n631), .B1(new_n581), .B2(new_n582), .ZN(new_n910));
  INV_X1    g485(.A(new_n582), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n632), .A3(new_n580), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n865), .B(new_n643), .Z(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n913), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT106), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n906), .A2(new_n909), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n906), .B2(new_n909), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n862), .A2(new_n635), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(G171), .A2(G286), .ZN(new_n934));
  NAND4_X1  g509(.A1(G301), .A2(new_n532), .A3(new_n534), .A4(new_n542), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n865), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n863), .A2(new_n934), .A3(new_n864), .A4(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n917), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT109), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n915), .B2(new_n916), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n913), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n939), .A2(new_n913), .A3(KEYINPUT110), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n942), .A2(new_n904), .A3(new_n945), .A4(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n951), .A2(new_n890), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n942), .A2(new_n945), .A3(new_n950), .ZN(new_n953));
  INV_X1    g528(.A(new_n904), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n933), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n890), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n946), .B1(new_n943), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n943), .A2(new_n958), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n904), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n957), .A2(new_n962), .A3(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n932), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT112), .B1(new_n957), .B2(new_n962), .ZN(new_n965));
  INV_X1    g540(.A(new_n961), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n954), .B1(new_n966), .B2(new_n959), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n951), .A3(new_n968), .A4(new_n890), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n965), .A2(KEYINPUT43), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n952), .A2(new_n933), .A3(new_n955), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n964), .B1(new_n970), .B2(new_n972), .ZN(G397));
  OAI21_X1  g548(.A(G40), .B1(new_n476), .B2(new_n463), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n474), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G164), .B2(G1384), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n739), .B(new_n741), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n718), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT127), .ZN(new_n983));
  INV_X1    g558(.A(G1996), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT46), .Z(new_n986));
  NOR2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  NOR2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n979), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(KEYINPUT48), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(KEYINPUT48), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n837), .A2(new_n839), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n717), .B(new_n984), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n837), .A2(new_n839), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n994), .A2(new_n981), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n992), .B(new_n993), .C1(new_n979), .C2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n837), .A2(new_n839), .A3(new_n981), .A4(new_n995), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n734), .A2(new_n738), .A3(new_n741), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n980), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n988), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1981), .B1(new_n545), .B2(G48), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n602), .A2(new_n606), .A3(new_n609), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n607), .B1(new_n519), .B2(new_n598), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n608), .A2(new_n504), .ZN(new_n1007));
  OAI21_X1  g582(.A(G1981), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT49), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G164), .A2(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n975), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1004), .A2(KEYINPUT49), .A3(new_n1008), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G288), .A2(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1005), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1012), .B(KEYINPUT117), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n813), .A2(new_n814), .A3(G1976), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1012), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1028), .A3(new_n1024), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1018), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  INV_X1    g606(.A(new_n502), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n501), .B1(new_n462), .B2(new_n498), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT45), .B(new_n1031), .C1(new_n1034), .C2(new_n496), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n978), .A2(new_n975), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1037));
  INV_X1    g612(.A(G1971), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n978), .A2(new_n975), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1043), .B(new_n1031), .C1(new_n1034), .C2(new_n496), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n975), .A3(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1045), .A2(G2090), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(G8), .B(new_n1049), .C1(new_n517), .C2(new_n523), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G166), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(new_n1055), .A3(G8), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1020), .A2(new_n1021), .B1(new_n1030), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1047), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1055), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1029), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1025), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1063), .A3(new_n1018), .A4(new_n1056), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT45), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(G164), .B2(G1384), .ZN(new_n1066));
  INV_X1    g641(.A(new_n977), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1031), .B(new_n1067), .C1(new_n1034), .C2(new_n496), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n975), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n730), .ZN(new_n1070));
  INV_X1    g645(.A(G2084), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1042), .A2(new_n975), .A3(new_n1044), .A4(new_n1071), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1051), .B(G286), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1058), .B1(new_n1064), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1056), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1055), .B1(new_n1047), .B2(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1030), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(KEYINPUT63), .A4(new_n1073), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1057), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1956), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1045), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n978), .A2(new_n975), .A3(new_n1035), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n573), .A2(new_n1087), .A3(new_n579), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n573), .B2(new_n579), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT119), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n573), .A2(new_n579), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT57), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n573), .A2(new_n1087), .A3(new_n579), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1086), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1086), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n631), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1045), .A2(new_n746), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n975), .A2(new_n1010), .A3(new_n741), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1097), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT122), .B1(new_n1086), .B2(new_n1098), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1109), .A2(new_n1096), .A3(KEYINPUT61), .A4(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT60), .B(new_n631), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1083), .A2(new_n1085), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1099), .B2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1011), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n978), .A2(new_n975), .A3(new_n1035), .A4(new_n984), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n559), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT121), .Z(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1121), .B(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT60), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT118), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1104), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1128), .A2(new_n1132), .A3(new_n632), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1108), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1061), .A2(new_n1056), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1070), .A2(G168), .A3(new_n1072), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G286), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(G8), .A3(new_n1136), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1141), .B2(KEYINPUT51), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1135), .A2(new_n1142), .A3(new_n1030), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1066), .A2(new_n975), .A3(new_n1068), .A4(new_n757), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1148));
  INV_X1    g723(.A(G1961), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1045), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(G2078), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1148), .B(new_n1150), .C1(KEYINPUT53), .C2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n1152), .B2(G171), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n757), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1155), .A2(new_n1144), .B1(new_n1149), .B2(new_n1045), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(G301), .A4(new_n1148), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n757), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1160));
  NAND4_X1  g735(.A1(G160), .A2(new_n978), .A3(new_n1035), .A4(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1150), .B(new_n1161), .C1(new_n1151), .C2(KEYINPUT53), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n1162), .B2(G171), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1153), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(G301), .B1(new_n1156), .B2(new_n1148), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(G171), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1134), .A2(new_n1143), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1081), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1081), .B2(new_n1168), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1141), .A2(KEYINPUT51), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1138), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1175), .A2(new_n1078), .A3(new_n1079), .A4(new_n1165), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1064), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1179), .A2(KEYINPUT126), .A3(new_n1165), .A4(new_n1175), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1142), .A2(new_n1173), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1170), .A2(new_n1171), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n997), .A2(new_n989), .ZN(new_n1184));
  NAND2_X1  g759(.A1(G290), .A2(G1986), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n980), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1002), .B1(new_n1183), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g762(.A1(new_n956), .A2(new_n963), .ZN(new_n1189));
  NOR3_X1   g763(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1190));
  OAI21_X1  g764(.A(new_n1190), .B1(new_n679), .B2(new_n678), .ZN(new_n1191));
  NOR3_X1   g765(.A1(new_n1189), .A2(new_n893), .A3(new_n1191), .ZN(G308));
  NOR2_X1   g766(.A1(new_n1191), .A2(new_n893), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(new_n956), .B2(new_n963), .ZN(G225));
endmodule


