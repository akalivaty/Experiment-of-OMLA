//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT65), .B(G77), .Z(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  AND3_X1   g0047(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(KEYINPUT25), .B1(new_n246), .B2(new_n247), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n245), .A2(new_n250), .A3(new_n216), .A4(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n248), .A2(new_n249), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT76), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT76), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n208), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n254), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G87), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(KEYINPUT22), .A3(G20), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n261), .A2(KEYINPUT22), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT76), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT76), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G116), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT23), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(new_n208), .B2(G107), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n247), .A2(KEYINPUT23), .A3(G20), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n276), .A2(new_n208), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT24), .B1(new_n271), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT24), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT22), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT3), .B1(new_n272), .B2(new_n273), .ZN(new_n285));
  AOI21_X1  g0085(.A(G20), .B1(new_n285), .B2(new_n265), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n286), .B2(G87), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n268), .A2(new_n270), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n283), .B(new_n280), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n251), .A2(new_n216), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n253), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT76), .B(G33), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n260), .B1(new_n293), .B2(KEYINPUT3), .ZN(new_n294));
  INV_X1    g0094(.A(G257), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G1698), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G250), .B2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G294), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n294), .A2(new_n297), .B1(new_n298), .B2(new_n274), .ZN(new_n299));
  AND2_X1   g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT68), .B1(new_n300), .B2(new_n216), .ZN(new_n301));
  AND2_X1   g0101(.A1(G1), .A2(G13), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n302), .B2(new_n304), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n207), .A2(G45), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT5), .B(G41), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n300), .A2(new_n216), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n311), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G264), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G190), .B2(new_n317), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n292), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G179), .B2(new_n317), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n292), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G20), .A2(G33), .ZN(new_n330));
  XOR2_X1   g0130(.A(new_n330), .B(KEYINPUT70), .Z(new_n331));
  NOR2_X1   g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n208), .A2(G33), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n219), .A2(new_n208), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n291), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n245), .A2(new_n216), .A3(new_n251), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n208), .A2(G1), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n337), .A2(new_n340), .B1(new_n219), .B2(new_n246), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT66), .ZN(new_n343));
  INV_X1    g0143(.A(G41), .ZN(new_n344));
  INV_X1    g0144(.A(G45), .ZN(new_n345));
  AOI21_X1  g0145(.A(G1), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n309), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n309), .B2(new_n346), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n314), .A2(new_n346), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n348), .A2(new_n349), .B1(new_n220), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n268), .A2(G232), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n268), .A2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G238), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n353), .B1(new_n247), .B2(new_n268), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n351), .B1(new_n356), .B2(new_n306), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n342), .B1(new_n357), .B2(G169), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(KEYINPUT71), .B1(new_n359), .B2(new_n357), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT71), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n342), .C1(new_n357), .C2(G169), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(G190), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n357), .A2(new_n318), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n342), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n360), .A2(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n368));
  INV_X1    g0168(.A(new_n291), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n327), .A2(new_n334), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(G150), .B2(new_n330), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n204), .A2(G20), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n338), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n337), .A2(G50), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G50), .B2(new_n245), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G223), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n354), .A2(new_n378), .B1(new_n219), .B2(new_n268), .ZN(new_n379));
  AOI21_X1  g0179(.A(G1698), .B1(new_n264), .B2(new_n267), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n380), .A2(G222), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n306), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n309), .A2(new_n346), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT66), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n314), .A2(new_n346), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n347), .B1(G226), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n377), .B1(new_n388), .B2(G169), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(G179), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT9), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n377), .A2(new_n393), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n373), .A2(new_n393), .A3(new_n376), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT10), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n394), .A2(new_n395), .ZN(new_n400));
  INV_X1    g0200(.A(new_n398), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .A4(new_n392), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n391), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n367), .A2(new_n368), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n337), .A2(G68), .A3(new_n374), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT74), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT75), .ZN(new_n408));
  AOI211_X1 g0208(.A(G68), .B(new_n245), .C1(new_n408), .C2(KEYINPUT12), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(KEYINPUT12), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n330), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n339), .B2(new_n334), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n291), .ZN(new_n415));
  XOR2_X1   g0215(.A(new_n415), .B(KEYINPUT11), .Z(new_n416));
  NOR2_X1   g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n355), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n380), .A2(G226), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n419), .B1(new_n423), .B2(new_n306), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n301), .A2(new_n305), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n380), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT73), .B1(new_n429), .B2(new_n419), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n426), .A2(new_n430), .A3(KEYINPUT13), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n359), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n424), .A2(new_n432), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n429), .B2(new_n419), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n322), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n434), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n435), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n418), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n378), .A2(new_n352), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G226), .B2(new_n352), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n294), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n256), .A2(new_n269), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n306), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n384), .A2(new_n347), .B1(G232), .B2(new_n385), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n447), .A2(G179), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n322), .B1(new_n447), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(G58), .B(G68), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(G20), .B1(G159), .B2(new_n330), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT7), .ZN(new_n454));
  NOR4_X1   g0254(.A1(new_n259), .A2(new_n454), .A3(G20), .A4(new_n260), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT77), .B1(new_n259), .B2(new_n260), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n285), .A2(new_n457), .A3(new_n265), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n208), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT16), .B(new_n453), .C1(new_n460), .C2(new_n203), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n264), .A2(new_n267), .A3(new_n208), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n274), .A2(new_n254), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n263), .A2(new_n454), .A3(G20), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n462), .A2(new_n454), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n453), .B1(new_n465), .B2(new_n203), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT16), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n369), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n327), .A2(new_n338), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n470), .A2(new_n337), .B1(new_n246), .B2(new_n327), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n451), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT18), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n447), .A2(new_n397), .A3(new_n448), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n447), .A2(new_n448), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(G200), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n476), .A3(new_n471), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT17), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n471), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n461), .B2(new_n468), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT17), .A3(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n431), .A2(G190), .A3(new_n436), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n424), .A2(new_n432), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n429), .A2(KEYINPUT13), .A3(new_n419), .ZN(new_n487));
  OAI21_X1  g0287(.A(G200), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n488), .A3(new_n417), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n442), .A2(new_n473), .A3(new_n484), .A4(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n405), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n462), .A2(new_n454), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n463), .A2(new_n464), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT78), .A3(G107), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT78), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n465), .B2(new_n247), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n247), .A2(KEYINPUT6), .A3(G97), .ZN(new_n498));
  XOR2_X1   g0298(.A(G97), .B(G107), .Z(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n330), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n291), .ZN(new_n503));
  INV_X1    g0303(.A(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n246), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n252), .B2(new_n504), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n315), .A2(G257), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n313), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n352), .A2(G244), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n294), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n511), .A2(new_n220), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n263), .A2(new_n260), .A3(new_n262), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT67), .B1(new_n265), .B2(new_n266), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n352), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  AOI211_X1 g0320(.A(G179), .B(new_n510), .C1(new_n520), .C2(new_n306), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n514), .A2(new_n519), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n512), .B1(new_n285), .B2(new_n265), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n515), .B1(new_n523), .B2(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n306), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n510), .ZN(new_n526));
  AOI21_X1  g0326(.A(G169), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n508), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n506), .B1(new_n502), .B2(new_n291), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n526), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G190), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n510), .B1(new_n520), .B2(new_n306), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT21), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n515), .B(new_n208), .C1(G33), .C2(new_n504), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n275), .A2(G20), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n291), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT20), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n246), .A2(new_n275), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n252), .B2(new_n275), .ZN(new_n547));
  OAI21_X1  g0347(.A(G169), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n312), .A2(new_n311), .ZN(new_n549));
  INV_X1    g0349(.A(new_n314), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(G270), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n313), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n352), .A2(G264), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n295), .A2(new_n352), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G303), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n294), .A2(new_n555), .B1(new_n268), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n552), .B1(new_n557), .B2(new_n306), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n537), .B1(new_n548), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(G190), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n545), .A2(new_n547), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n318), .C2(new_n558), .ZN(new_n562));
  INV_X1    g0362(.A(new_n558), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n544), .B(new_n546), .C1(new_n275), .C2(new_n252), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT21), .A4(G169), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n359), .B(new_n552), .C1(new_n306), .C2(new_n557), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n564), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n559), .A2(new_n562), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n355), .A2(new_n352), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n220), .A2(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n285), .B2(new_n265), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n306), .B1(new_n573), .B2(new_n276), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n310), .A2(G250), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n550), .A2(new_n575), .B1(new_n309), .B2(new_n311), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n574), .A2(G179), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n322), .B1(new_n574), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(G179), .A3(new_n576), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n259), .B2(new_n260), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n293), .A2(G116), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n427), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n576), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(KEYINPUT79), .B(new_n580), .C1(new_n586), .C2(new_n322), .ZN(new_n587));
  INV_X1    g0387(.A(new_n333), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n245), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT80), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n337), .A2(new_n588), .A3(new_n591), .A4(new_n250), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT80), .B1(new_n252), .B2(new_n333), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(G20), .B1(G33), .B2(G97), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT19), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OR3_X1    g0397(.A1(new_n334), .A2(KEYINPUT19), .A3(new_n504), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n286), .A2(G68), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n590), .B(new_n594), .C1(new_n599), .C2(new_n369), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n579), .A2(new_n587), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n584), .B2(new_n585), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n208), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n598), .A2(new_n597), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n589), .B1(new_n605), .B2(new_n291), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n252), .A2(new_n269), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT81), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n574), .A2(G190), .A3(new_n576), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n602), .A2(new_n606), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n568), .A2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n326), .A2(new_n491), .A3(new_n536), .A4(new_n613), .ZN(G372));
  NAND3_X1  g0414(.A1(new_n489), .A2(new_n362), .A3(new_n360), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n483), .B1(new_n442), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT18), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n472), .B(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n399), .B2(new_n403), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(new_n391), .ZN(new_n621));
  INV_X1    g0421(.A(new_n491), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT26), .B1(new_n529), .B2(new_n612), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n530), .A2(new_n521), .A3(new_n527), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n600), .B1(new_n577), .B2(new_n578), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n611), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n623), .A2(new_n629), .A3(new_n626), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n292), .B2(new_n320), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT82), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n631), .A2(new_n529), .A3(new_n535), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n559), .A2(new_n565), .A3(new_n567), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n292), .A2(new_n324), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n631), .A2(new_n529), .A3(new_n535), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT82), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n630), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n621), .B1(new_n622), .B2(new_n641), .ZN(G369));
  INV_X1    g0442(.A(KEYINPUT83), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n561), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n643), .B1(new_n568), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n634), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n634), .A2(new_n643), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT84), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT84), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(new_n658), .A3(new_n655), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(G330), .A3(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT86), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n636), .B2(new_n650), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n325), .A2(KEYINPUT86), .A3(new_n649), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n292), .A2(new_n650), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n326), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n635), .A2(new_n649), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n636), .A2(new_n649), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n211), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n595), .A2(new_n275), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n680), .A2(new_n207), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n215), .ZN(new_n683));
  INV_X1    g0483(.A(new_n680), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n682), .A2(KEYINPUT87), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(KEYINPUT87), .B2(new_n682), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT28), .Z(new_n687));
  NAND3_X1  g0487(.A1(new_n640), .A2(new_n637), .A3(new_n633), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n623), .A2(new_n629), .A3(new_n626), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n649), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT89), .B1(new_n690), .B2(KEYINPUT29), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n692), .B(new_n693), .C1(new_n641), .C2(new_n649), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n529), .B2(new_n627), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n626), .B(KEYINPUT90), .Z(new_n696));
  NAND3_X1  g0496(.A1(new_n624), .A2(new_n611), .A3(new_n601), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(KEYINPUT26), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n639), .B1(new_n636), .B2(new_n635), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT29), .B(new_n650), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n691), .A2(new_n694), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n299), .A2(new_n306), .B1(new_n315), .B2(G264), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n558), .A2(new_n586), .A3(new_n704), .A4(G179), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT88), .B(new_n703), .C1(new_n705), .C2(new_n531), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n558), .A2(new_n586), .A3(G179), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(new_n317), .A3(new_n531), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n586), .A2(new_n704), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(KEYINPUT88), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n566), .A3(new_n533), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n706), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n712), .B2(new_n649), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n536), .A2(new_n326), .A3(new_n613), .A4(new_n650), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n702), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n687), .B1(new_n720), .B2(G1), .ZN(G364));
  AND2_X1   g0521(.A1(new_n208), .A2(G13), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n207), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n680), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(G330), .B1(new_n657), .B2(new_n659), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n663), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n657), .B2(new_n659), .ZN(new_n733));
  INV_X1    g0533(.A(new_n268), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n679), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G355), .B1(new_n275), .B2(new_n679), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n243), .A2(G45), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G45), .B2(new_n683), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n456), .A2(new_n458), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n679), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n736), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n216), .B1(G20), .B2(new_n322), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n731), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n397), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n359), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n208), .A2(new_n359), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n749), .A2(new_n298), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n397), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(KEYINPUT92), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(KEYINPUT92), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n754), .B1(new_n760), .B2(G326), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT95), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n208), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n734), .B1(new_n556), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(KEYINPUT96), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT96), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n755), .A2(G190), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n763), .A2(new_n751), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n768), .A2(new_n769), .B1(G329), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n750), .A2(new_n746), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT91), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(KEYINPUT91), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n767), .B(new_n772), .C1(new_n773), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n763), .A2(new_n397), .A3(G200), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT93), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n766), .B(new_n779), .C1(G283), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(G107), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n748), .A2(G97), .ZN(new_n789));
  OAI21_X1  g0589(.A(KEYINPUT32), .B1(new_n770), .B2(new_n787), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n219), .ZN(new_n792));
  INV_X1    g0592(.A(new_n752), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n734), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n764), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n768), .A2(G68), .B1(new_n795), .B2(G87), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(new_n202), .C2(new_n778), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n791), .B(new_n797), .C1(G50), .C2(new_n760), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n762), .A2(new_n785), .B1(new_n786), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n743), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n745), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n725), .B1(new_n733), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n728), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT97), .Z(G396));
  NAND2_X1  g0604(.A1(new_n688), .A2(new_n689), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n366), .A2(new_n650), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT99), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT99), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n809), .B(new_n806), .C1(new_n688), .C2(new_n689), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n357), .A2(new_n359), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n811), .A2(new_n362), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n365), .A2(new_n363), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n650), .B1(new_n336), .B2(new_n341), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n813), .B2(new_n816), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n808), .A2(new_n810), .B1(new_n690), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n725), .B1(new_n819), .B2(new_n718), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n718), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n743), .A2(new_n729), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT98), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n725), .B1(new_n823), .B2(G77), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n734), .B1(new_n275), .B2(new_n752), .C1(new_n753), .C2(new_n770), .ZN(new_n825));
  INV_X1    g0625(.A(new_n768), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n789), .B1(new_n247), .B2(new_n764), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n778), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n825), .B(new_n828), .C1(G294), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n784), .A2(G87), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(new_n556), .C2(new_n759), .ZN(new_n832));
  INV_X1    g0632(.A(new_n739), .ZN(new_n833));
  INV_X1    g0633(.A(new_n784), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n203), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n749), .A2(new_n202), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n764), .A2(new_n201), .B1(new_n770), .B2(new_n837), .ZN(new_n838));
  OR4_X1    g0638(.A1(new_n833), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n768), .A2(G150), .B1(new_n793), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n841), .B2(new_n778), .C1(new_n759), .C2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  OAI21_X1  g0644(.A(new_n832), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n824), .B1(new_n845), .B2(new_n743), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n818), .B2(new_n730), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n821), .A2(KEYINPUT100), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT100), .B1(new_n821), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  OR2_X1    g0651(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(G116), .A3(new_n217), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT36), .Z(new_n855));
  OAI211_X1 g0655(.A(new_n215), .B(new_n792), .C1(new_n202), .C2(new_n203), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n203), .A2(G50), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT101), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n207), .B(G13), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n360), .A2(new_n362), .A3(new_n650), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n808), .B2(new_n810), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n453), .B1(new_n460), .B2(new_n203), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n467), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n461), .A2(new_n291), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n471), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n451), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n647), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n871), .A3(new_n477), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n477), .B1(new_n481), .B2(new_n451), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n481), .B2(new_n647), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n469), .A2(new_n471), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n868), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(KEYINPUT103), .A3(new_n880), .A4(new_n477), .ZN(new_n881));
  AOI22_X1  g0681(.A1(KEYINPUT37), .A2(new_n872), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n871), .B1(new_n473), .B2(new_n484), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n863), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n877), .A2(new_n881), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n870), .B(new_n867), .C1(new_n618), .C2(new_n483), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(G169), .B1(new_n486), .B2(new_n487), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(KEYINPUT14), .B1(new_n431), .B2(new_n433), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n417), .B1(new_n892), .B2(new_n440), .ZN(new_n893));
  INV_X1    g0693(.A(new_n489), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n418), .B2(new_n649), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n417), .A2(KEYINPUT102), .A3(new_n650), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n893), .A2(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n442), .A2(new_n489), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n862), .A2(new_n890), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n618), .A2(new_n647), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n481), .A2(new_n647), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n618), .B2(new_n483), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n877), .A2(new_n881), .A3(KEYINPUT106), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n874), .B2(new_n904), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT106), .B1(new_n877), .B2(new_n881), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n882), .A2(new_n883), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT39), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n915), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT104), .B1(new_n442), .B2(new_n649), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT104), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n893), .A2(new_n918), .A3(new_n650), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n902), .B(new_n903), .C1(new_n916), .C2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n621), .B1(new_n701), .B2(new_n622), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n882), .A2(new_n863), .A3(new_n883), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n887), .B2(new_n888), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n715), .A2(new_n716), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n929), .A2(new_n818), .A3(new_n898), .A4(new_n900), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n925), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n925), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n886), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n907), .A3(new_n906), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n911), .B1(new_n935), .B2(new_n905), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n932), .B1(new_n936), .B2(new_n926), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n491), .A2(new_n929), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(G330), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n924), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n207), .B2(new_n722), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n924), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n860), .B1(new_n944), .B2(new_n945), .ZN(G367));
  OAI21_X1  g0746(.A(new_n536), .B1(new_n530), .B2(new_n650), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n624), .A2(new_n649), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n673), .A2(new_n950), .A3(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT42), .B1(new_n673), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n529), .B1(new_n947), .B2(new_n636), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n650), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n606), .A2(new_n609), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n649), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(new_n626), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT107), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n959), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n960), .B(new_n961), .C1(new_n627), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT43), .Z(new_n966));
  AND3_X1   g0766(.A1(new_n956), .A2(new_n957), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n965), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n956), .B2(new_n957), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n671), .A2(new_n950), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n967), .A2(new_n970), .B1(new_n971), .B2(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT109), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n680), .B(KEYINPUT41), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n676), .A2(new_n950), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT110), .B1(new_n677), .B2(new_n949), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT110), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n676), .A2(new_n980), .A3(new_n950), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n981), .A3(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT44), .B1(new_n979), .B2(new_n981), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n663), .B(new_n670), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT111), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n670), .A2(new_n672), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n673), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n663), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n661), .A2(new_n662), .A3(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n986), .B1(new_n992), .B2(new_n719), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n661), .A2(new_n662), .A3(new_n988), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n988), .B1(new_n661), .B2(new_n662), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(KEYINPUT111), .A3(new_n720), .ZN(new_n997));
  INV_X1    g0797(.A(new_n984), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n998), .A2(new_n671), .A3(new_n978), .A4(new_n982), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n985), .A2(new_n993), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n976), .B1(new_n1000), .B2(new_n720), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n974), .B(new_n975), .C1(new_n1001), .C2(new_n724), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n744), .B1(new_n211), .B2(new_n333), .C1(new_n741), .C2(new_n236), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(new_n725), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n759), .A2(new_n753), .B1(new_n504), .B2(new_n783), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n752), .A2(new_n827), .B1(new_n770), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G107), .B2(new_n748), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n833), .C1(new_n298), .C2(new_n826), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT46), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n764), .B2(new_n275), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n778), .C2(new_n556), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1005), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n748), .A2(G68), .ZN(new_n1015));
  INV_X1    g0815(.A(G150), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n1016), .B2(new_n778), .C1(new_n759), .C2(new_n841), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT112), .Z(new_n1018));
  AOI22_X1  g0818(.A1(new_n768), .A2(G159), .B1(new_n795), .B2(G58), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G50), .A2(new_n793), .B1(new_n771), .B2(G137), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n268), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n783), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1021), .B1(new_n792), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1014), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1004), .B1(new_n732), .B2(new_n968), .C1(new_n1025), .C2(new_n800), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1002), .A2(new_n1026), .ZN(G387));
  NAND2_X1  g0827(.A1(new_n993), .A2(new_n997), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n684), .B1(new_n992), .B2(new_n719), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n996), .A2(new_n724), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n826), .A2(new_n327), .B1(new_n749), .B2(new_n333), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G68), .A2(new_n793), .B1(new_n771), .B2(G150), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n219), .B2(new_n764), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G50), .C2(new_n829), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n833), .B1(new_n760), .B2(G159), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n504), .C2(new_n834), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n739), .B1(G326), .B2(new_n771), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n749), .A2(new_n827), .B1(new_n764), .B2(new_n298), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n768), .A2(G311), .B1(new_n793), .B2(G303), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n1006), .B2(new_n778), .C1(new_n759), .C2(new_n773), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1038), .B1(new_n275), .B2(new_n783), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1037), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n743), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n735), .A2(new_n681), .B1(new_n247), .B2(new_n679), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n329), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n201), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n345), .B1(new_n203), .B2(new_n339), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1053), .A2(new_n681), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n740), .B1(new_n233), .B2(new_n345), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n726), .B1(new_n1057), .B2(new_n744), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1049), .B(new_n1058), .C1(new_n670), .C2(new_n732), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1030), .A2(new_n1031), .A3(new_n1059), .ZN(G393));
  AND2_X1   g0860(.A1(new_n985), .A2(new_n999), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n724), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n744), .B1(new_n504), .B2(new_n211), .C1(new_n741), .C2(new_n240), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n725), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n759), .A2(new_n1006), .B1(new_n753), .B2(new_n778), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT52), .Z(new_n1066));
  AOI22_X1  g0866(.A1(G116), .A2(new_n748), .B1(new_n793), .B2(G294), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n556), .B2(new_n826), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n770), .A2(new_n773), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1070), .B(new_n268), .C1(G283), .C2(new_n795), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n786), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n759), .A2(new_n1016), .B1(new_n787), .B2(new_n778), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  AOI22_X1  g0874(.A1(new_n768), .A2(G50), .B1(new_n795), .B2(G68), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n748), .A2(G77), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n841), .C2(new_n770), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1051), .B2(new_n793), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n831), .A2(new_n1078), .A3(new_n739), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1066), .A2(new_n1072), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1064), .B1(new_n1080), .B2(new_n743), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n949), .B2(new_n732), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1000), .A2(new_n680), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n999), .A2(new_n985), .B1(new_n993), .B2(new_n997), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1062), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(G390));
  NAND2_X1  g0885(.A1(new_n916), .A2(new_n729), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n823), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1087), .A2(new_n327), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n734), .B1(new_n504), .B2(new_n752), .C1(new_n298), .C2(new_n770), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1076), .B1(new_n269), .B2(new_n764), .C1(new_n826), .C2(new_n247), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G116), .C2(new_n829), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n827), .B2(new_n759), .ZN(new_n1092));
  OR3_X1    g0892(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n1016), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT53), .B1(new_n764), .B2(new_n1016), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n778), .C2(new_n837), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n760), .A2(G128), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n826), .A2(new_n842), .B1(new_n749), .B2(new_n787), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  INV_X1    g0898(.A(G125), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n752), .A2(new_n1098), .B1(new_n770), .B2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1097), .A2(new_n734), .A3(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1096), .B(new_n1101), .C1(new_n201), .C2(new_n783), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1092), .A2(new_n835), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n800), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n726), .B(new_n1088), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1086), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n818), .B(new_n650), .C1(new_n698), .C2(new_n699), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n861), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n920), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n917), .A2(KEYINPUT114), .A3(new_n919), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1110), .A2(new_n901), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n926), .B2(new_n936), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n920), .B1(new_n862), .B2(new_n901), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT39), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n889), .A2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n928), .A2(new_n1117), .B1(new_n936), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n717), .A2(new_n818), .A3(new_n900), .A4(new_n898), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1115), .B(new_n1121), .C1(new_n1116), .C2(new_n1119), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1108), .B1(new_n1125), .B2(new_n723), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n929), .A2(G330), .A3(new_n818), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n898), .A2(new_n900), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1121), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n862), .A2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1109), .A2(new_n861), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n1130), .A3(new_n1121), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n491), .A2(new_n717), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n621), .B(new_n1136), .C1(new_n701), .C2(new_n622), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n684), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1123), .A2(new_n1124), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT115), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1124), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n861), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n809), .B1(new_n641), .B2(new_n806), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n805), .A2(KEYINPUT99), .A3(new_n807), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n921), .B1(new_n1147), .B2(new_n1129), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n916), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1121), .B1(new_n1149), .B2(new_n1115), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1138), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  AND4_X1   g0951(.A1(KEYINPUT115), .A2(new_n1151), .A3(new_n680), .A4(new_n1141), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1127), .B1(new_n1142), .B2(new_n1152), .ZN(G378));
  NAND2_X1  g0953(.A1(new_n377), .A2(new_n870), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT55), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n404), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n404), .A2(new_n1157), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1160), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1156), .B(new_n391), .C1(new_n399), .C2(new_n403), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n930), .B1(new_n884), .B2(new_n889), .ZN(new_n1167));
  OAI21_X1  g0967(.A(G330), .B1(new_n1167), .B2(KEYINPUT40), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n929), .A4(new_n818), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n913), .B2(new_n889), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1166), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT119), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1160), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1158), .A2(new_n1164), .A3(new_n1163), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1162), .A2(new_n1165), .A3(KEYINPUT119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n931), .A2(new_n937), .A3(new_n1177), .A4(G330), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n916), .A2(new_n921), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n902), .A2(new_n903), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n922), .A2(new_n1171), .A3(new_n1178), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n724), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n726), .B1(new_n201), .B2(new_n822), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n764), .A2(new_n1098), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT117), .Z(new_n1188));
  AOI22_X1  g0988(.A1(G150), .A2(new_n748), .B1(new_n793), .B2(G137), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n837), .B2(new_n826), .C1(new_n759), .C2(new_n1099), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(G128), .C2(new_n829), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT59), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1022), .A2(G159), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G33), .B(G41), .C1(new_n771), .C2(G124), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1022), .A2(G58), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n833), .C1(new_n275), .C2(new_n759), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1015), .B1(new_n219), .B2(new_n764), .C1(new_n826), .C2(new_n504), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n778), .A2(new_n247), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n344), .B1(new_n770), .B2(new_n827), .C1(new_n333), .C2(new_n752), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n344), .B1(new_n833), .B2(new_n256), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n201), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1197), .A2(new_n1204), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1186), .B1(new_n800), .B2(new_n1208), .C1(new_n1177), .C2(new_n730), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1185), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1137), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1141), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n680), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1141), .A2(new_n1212), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n922), .A2(new_n1171), .A3(new_n1178), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n922), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1211), .B1(new_n1215), .B2(new_n1220), .ZN(G375));
  NAND2_X1  g1021(.A1(new_n760), .A2(G294), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n764), .A2(new_n504), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n749), .A2(new_n333), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G116), .C2(new_n768), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n829), .A2(G283), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n752), .A2(new_n247), .B1(new_n770), .B2(new_n556), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(new_n268), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1222), .A2(new_n1225), .A3(new_n1226), .A4(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n834), .A2(new_n339), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G150), .A2(new_n793), .B1(new_n771), .B2(G128), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n826), .B2(new_n1098), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n795), .A2(G159), .B1(new_n748), .B2(G50), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n842), .C2(new_n778), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1198), .B(new_n739), .C1(new_n837), .C2(new_n759), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1229), .A2(new_n1230), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n743), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n726), .B1(new_n1087), .B2(new_n203), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n901), .C2(new_n730), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1135), .B2(new_n723), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT120), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n976), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1138), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(G381));
  NOR3_X1   g1046(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT121), .Z(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1126), .B1(new_n1141), .B2(new_n1139), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1242), .A3(new_n1245), .A4(new_n1250), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G387), .A2(new_n1248), .A3(G375), .A4(new_n1251), .ZN(G407));
  NAND2_X1  g1052(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT57), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n684), .B1(new_n1256), .B2(new_n1216), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1210), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n648), .A2(G213), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT122), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1250), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G407), .A2(G213), .A3(new_n1261), .ZN(G409));
  OAI21_X1  g1062(.A(KEYINPUT123), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT123), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1183), .A2(new_n1264), .A3(new_n1184), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n724), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1216), .A2(new_n1219), .A3(new_n1243), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1209), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1250), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1151), .A2(new_n680), .A3(new_n1141), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT115), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1139), .A2(KEYINPUT115), .A3(new_n1141), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1126), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1269), .B1(G375), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1260), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1140), .A2(new_n684), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1244), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1244), .A2(KEYINPUT124), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1242), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n850), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1279), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1277), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G384), .A3(new_n1242), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1275), .A2(new_n1276), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1260), .A2(G2897), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1285), .A2(new_n1288), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1290), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  XOR2_X1   g1098(.A(G393), .B(G396), .Z(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1002), .A2(new_n1026), .A3(G390), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G390), .B1(new_n1002), .B2(new_n1026), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(new_n1249), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1002), .A2(new_n1026), .A3(G390), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1299), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1303), .A2(new_n1306), .A3(KEYINPUT125), .A4(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1258), .A2(G378), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1260), .B1(new_n1312), .B2(new_n1269), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1298), .A2(new_n1308), .A3(new_n1311), .A4(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1275), .A2(new_n1276), .A3(new_n1289), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1313), .B2(new_n1289), .ZN(new_n1322));
  OAI211_X1 g1122(.A(KEYINPUT127), .B(new_n1316), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1290), .A2(new_n1317), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(new_n1320), .A3(new_n1319), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1327), .B2(new_n1316), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1315), .B1(new_n1325), .B2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1250), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1330), .A2(new_n1312), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1289), .ZN(new_n1332));
  XOR2_X1   g1132(.A(new_n1332), .B(new_n1324), .Z(G402));
endmodule


