//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT69), .A2(G953), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT69), .A2(G953), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n194), .A3(G214), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n194), .A3(G143), .A4(G214), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT18), .A2(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n201), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n198), .A3(new_n203), .A4(new_n199), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT75), .A2(G140), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT75), .A2(G140), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT76), .B(G125), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  OR2_X1    g023(.A1(KEYINPUT75), .A2(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT75), .A2(G140), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(G140), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n208), .B(G146), .C1(new_n212), .C2(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n209), .A2(G140), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n213), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT69), .B(G953), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT68), .B(G237), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(G143), .B1(new_n224), .B2(G214), .ZN(new_n225));
  INV_X1    g039(.A(new_n199), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n197), .A2(new_n228), .A3(new_n199), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n208), .B(KEYINPUT16), .C1(new_n212), .C2(new_n215), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT16), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n208), .B(KEYINPUT19), .C1(new_n212), .C2(new_n215), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT19), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n217), .A2(new_n213), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n218), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G113), .B(G122), .ZN(new_n242));
  INV_X1    g056(.A(G104), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n221), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(G475), .A2(G902), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n202), .A2(new_n204), .B1(new_n219), .B2(new_n216), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT17), .B(G131), .C1(new_n225), .C2(new_n226), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n231), .A2(new_n218), .A3(new_n233), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(new_n250), .A3(new_n235), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n227), .A2(new_n252), .A3(new_n229), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n246), .B(new_n247), .C1(new_n254), .C2(new_n245), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT20), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n257));
  INV_X1    g071(.A(new_n247), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT87), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n259), .B2(new_n258), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n246), .B(new_n261), .C1(new_n254), .C2(new_n245), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT88), .ZN(new_n263));
  INV_X1    g077(.A(new_n250), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n218), .B1(new_n231), .B2(new_n233), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n253), .A2(new_n266), .A3(new_n249), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n244), .B1(new_n267), .B2(new_n248), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n269), .A3(new_n246), .A4(new_n261), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n256), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT94), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT74), .B(G902), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G143), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n196), .A2(G128), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n196), .A2(G128), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT13), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n275), .A2(KEYINPUT93), .A3(KEYINPUT13), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n278), .B2(new_n279), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n277), .B1(new_n284), .B2(G134), .ZN(new_n285));
  INV_X1    g099(.A(G107), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT91), .A2(G122), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(KEYINPUT91), .A2(G122), .ZN(new_n289));
  OAI21_X1  g103(.A(G116), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT91), .B(G122), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT92), .A3(G116), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G116), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G122), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n286), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  AOI211_X1 g113(.A(G107), .B(new_n299), .C1(new_n292), .C2(new_n294), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n285), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n286), .A3(new_n297), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n275), .A2(new_n276), .ZN(new_n303));
  INV_X1    g117(.A(G134), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n297), .B(KEYINPUT14), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n292), .B2(new_n294), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n302), .B(new_n305), .C1(new_n286), .C2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(new_n310), .A3(G953), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n301), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n301), .B2(new_n308), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n272), .B(new_n273), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G478), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT15), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n314), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n312), .ZN(new_n320));
  INV_X1    g134(.A(new_n317), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n272), .A3(new_n273), .A4(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(G952), .ZN(new_n325));
  NAND2_X1  g139(.A1(G234), .A2(G237), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n327), .B(KEYINPUT95), .Z(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n273), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n326), .A3(new_n222), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT21), .B(G898), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n244), .A2(KEYINPUT90), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n267), .B2(new_n248), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n251), .A2(new_n253), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n336), .A3(new_n221), .ZN(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT89), .B(G475), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n271), .A2(new_n323), .A3(new_n335), .A4(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT96), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n218), .A2(G143), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n196), .A2(G146), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G143), .B2(new_n218), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n351), .B2(new_n274), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n347), .A2(new_n348), .A3(new_n350), .A4(G128), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n209), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n324), .A2(G224), .ZN(new_n356));
  NOR2_X1   g170(.A1(KEYINPUT0), .A2(G128), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(KEYINPUT0), .A2(G128), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n349), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G143), .B(G146), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n359), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n355), .B(new_n356), .C1(new_n209), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n357), .B1(new_n362), .B2(new_n359), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n349), .A2(new_n360), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n209), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G125), .B1(new_n352), .B2(new_n353), .ZN(new_n369));
  OAI211_X1 g183(.A(G224), .B(new_n324), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n286), .A3(KEYINPUT3), .A4(G104), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n243), .A2(KEYINPUT81), .A3(G107), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n286), .B2(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n374), .C1(new_n375), .C2(new_n377), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n243), .A2(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n286), .A2(G104), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n376), .B(new_n384), .C1(new_n385), .C2(KEYINPUT81), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n381), .B1(new_n386), .B2(new_n374), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n380), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n378), .A2(KEYINPUT82), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n372), .A3(G101), .A4(new_n382), .ZN(new_n390));
  XNOR2_X1  g204(.A(G116), .B(G119), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(KEYINPUT2), .A2(G113), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT66), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(KEYINPUT2), .B2(G113), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT2), .A2(G113), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT67), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n392), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n394), .A2(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n391), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(new_n390), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n379), .B1(new_n385), .B2(new_n384), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n378), .B2(new_n379), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G116), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(G113), .C1(KEYINPUT5), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n413), .A3(new_n405), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G122), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n407), .A2(new_n414), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n416), .A2(KEYINPUT6), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n371), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT7), .B1(new_n324), .B2(G224), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n365), .A2(new_n370), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n378), .A2(new_n379), .ZN(new_n426));
  INV_X1    g240(.A(new_n408), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n405), .A3(new_n413), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n415), .B(KEYINPUT8), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n410), .A2(KEYINPUT85), .ZN(new_n431));
  OAI21_X1  g245(.A(G113), .B1(new_n412), .B2(KEYINPUT5), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n410), .B2(KEYINPUT85), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n431), .A2(new_n433), .B1(new_n391), .B2(new_n404), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n429), .B(new_n430), .C1(new_n434), .C2(new_n428), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n355), .B(new_n423), .C1(new_n209), .C2(new_n364), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n425), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n437), .B2(new_n416), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n422), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G210), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n422), .A2(new_n438), .A3(new_n440), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n346), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n310), .B1(new_n273), .B2(G234), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT23), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n411), .B2(G128), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n411), .A2(G128), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n274), .A2(KEYINPUT23), .A3(G119), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT77), .ZN(new_n458));
  INV_X1    g272(.A(G110), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n274), .A2(G119), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n455), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT24), .B(G110), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT77), .B1(new_n465), .B2(G110), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n219), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n467), .A2(new_n265), .A3(new_n468), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n457), .A2(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n235), .B2(new_n250), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n452), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G137), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n470), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n264), .B2(new_n265), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n235), .A2(new_n478), .A3(new_n219), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT78), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n475), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT78), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT25), .B1(new_n484), .B2(new_n273), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n486), .B(new_n330), .C1(new_n481), .C2(new_n483), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n451), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n451), .A2(G902), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n488), .A2(KEYINPUT79), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT79), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G137), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G134), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(KEYINPUT65), .A2(G137), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT65), .A2(G137), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n496), .B1(new_n499), .B2(new_n304), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n354), .B1(new_n228), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT11), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n304), .B2(G137), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT64), .ZN(new_n504));
  AND2_X1   g318(.A1(KEYINPUT11), .A2(G134), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT64), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n495), .A2(new_n507), .A3(new_n502), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n494), .A2(G134), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n504), .A2(new_n506), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(G131), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n501), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(G131), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(new_n495), .B2(new_n502), .ZN(new_n515));
  AOI211_X1 g329(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n494), .C2(G134), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(KEYINPUT65), .A2(G137), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT65), .A2(G137), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n509), .B1(new_n520), .B2(new_n505), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n521), .A3(new_n228), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n364), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n513), .A2(new_n523), .A3(new_n406), .ZN(new_n524));
  INV_X1    g338(.A(new_n406), .ZN(new_n525));
  INV_X1    g339(.A(new_n364), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n228), .B1(new_n517), .B2(new_n521), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n512), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n522), .B(new_n354), .C1(new_n228), .C2(new_n500), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT28), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n224), .A2(G210), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT27), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n532), .B(KEYINPUT27), .ZN(new_n537));
  INV_X1    g351(.A(new_n535), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n541), .A2(KEYINPUT29), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n528), .A2(new_n525), .A3(new_n529), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(KEYINPUT70), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT70), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT72), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n524), .B2(KEYINPUT28), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n551), .B2(new_n545), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n531), .B(new_n542), .C1(new_n548), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  INV_X1    g368(.A(new_n531), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT72), .B1(new_n546), .B2(new_n547), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n549), .A3(new_n545), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n542), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n513), .A2(new_n523), .A3(KEYINPUT30), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n528), .B2(new_n529), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n406), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n543), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT29), .B1(new_n565), .B2(new_n540), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n531), .A2(new_n551), .A3(new_n545), .A4(new_n541), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n330), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n554), .A2(new_n560), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G472), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n543), .A3(new_n541), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT30), .B1(new_n513), .B2(new_n523), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n528), .A2(new_n562), .A3(new_n529), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n524), .B1(new_n576), .B2(new_n406), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT31), .A3(new_n541), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n531), .A2(new_n551), .A3(new_n545), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n573), .A2(new_n578), .B1(new_n579), .B2(new_n540), .ZN(new_n580));
  NOR2_X1   g394(.A1(G472), .A2(G902), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT71), .Z(new_n582));
  OAI21_X1  g396(.A(KEYINPUT32), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n540), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT31), .B1(new_n577), .B2(new_n541), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n525), .B1(new_n574), .B2(new_n575), .ZN(new_n586));
  NOR4_X1   g400(.A1(new_n586), .A2(new_n572), .A3(new_n540), .A4(new_n524), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  INV_X1    g403(.A(new_n582), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n570), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G469), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n341), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n194), .A2(G227), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT80), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n388), .A2(new_n526), .A3(new_n390), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n514), .A2(new_n522), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT10), .B1(new_n409), .B2(new_n354), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n409), .A2(KEYINPUT10), .A3(new_n354), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n603), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n409), .A2(KEYINPUT10), .A3(new_n354), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n606), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n605), .B1(new_n612), .B2(new_n603), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n602), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n409), .B(new_n354), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n615), .A2(KEYINPUT12), .A3(new_n604), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT12), .B1(new_n615), .B2(new_n604), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n609), .B(new_n601), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n330), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n597), .B1(new_n619), .B2(new_n596), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(new_n601), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT83), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT83), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n609), .A2(new_n623), .A3(new_n601), .ZN(new_n624));
  INV_X1    g438(.A(new_n613), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n609), .B1(new_n616), .B2(new_n617), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n602), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(G469), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n595), .B1(new_n620), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n493), .A2(new_n593), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n450), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT97), .B(G101), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G3));
  NAND2_X1  g448(.A1(new_n588), .A2(new_n273), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n588), .A2(new_n590), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n271), .A2(new_n344), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n320), .A2(new_n273), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n316), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT33), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n312), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n301), .A2(new_n308), .A3(KEYINPUT100), .A4(new_n311), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n301), .A2(new_n308), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT99), .ZN(new_n648));
  INV_X1    g462(.A(new_n311), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n301), .A2(new_n308), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n642), .B1(new_n653), .B2(KEYINPUT33), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n330), .A2(new_n316), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n641), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n639), .A2(new_n657), .A3(new_n335), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n442), .A2(KEYINPUT98), .A3(new_n444), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n422), .A2(new_n438), .A3(new_n660), .A4(new_n440), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n661), .A2(new_n447), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n493), .A2(new_n638), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT34), .B(G104), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  NAND4_X1  g481(.A1(new_n268), .A2(new_n257), .A3(new_n246), .A4(new_n247), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n256), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n318), .A2(new_n322), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n335), .A3(new_n670), .A4(new_n344), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n672), .A2(KEYINPUT101), .A3(new_n659), .A4(new_n662), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n663), .B2(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n493), .A3(new_n638), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NAND2_X1  g493(.A1(new_n477), .A2(new_n479), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT102), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n482), .A2(KEYINPUT36), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n489), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n488), .A2(new_n686), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n630), .A2(new_n636), .A3(new_n687), .A4(new_n637), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n346), .A2(new_n688), .A3(new_n449), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n329), .B1(new_n332), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n342), .B2(new_n343), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n669), .A2(new_n694), .A3(new_n670), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n687), .A2(new_n630), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n663), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n593), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XOR2_X1   g513(.A(new_n693), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n630), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT104), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n639), .A2(new_n670), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n687), .A3(new_n448), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n446), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n577), .A2(new_n540), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n524), .A2(new_n530), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n341), .B1(new_n710), .B2(new_n541), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n592), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n703), .A2(new_n704), .A3(new_n706), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n451), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n484), .A2(new_n273), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n486), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n484), .A2(KEYINPUT25), .A3(new_n273), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n684), .A2(new_n685), .A3(new_n489), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n630), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n693), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n639), .A2(new_n657), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n593), .A3(new_n697), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  OR2_X1    g543(.A1(new_n619), .A2(new_n596), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n619), .A2(new_n596), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n594), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n493), .A2(new_n593), .A3(new_n664), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n493), .A2(new_n593), .A3(new_n733), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n673), .A2(new_n675), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n569), .A2(G472), .B1(new_n583), .B2(new_n591), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n492), .A3(new_n491), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT105), .A3(new_n676), .A4(new_n733), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NOR2_X1   g559(.A1(new_n663), .A2(new_n732), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n346), .A2(new_n593), .A3(new_n687), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  OAI22_X1  g562(.A1(new_n558), .A2(new_n541), .B1(new_n585), .B2(new_n587), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n590), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n636), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n488), .A2(new_n490), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n705), .A2(new_n663), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n335), .A3(new_n733), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  AND3_X1   g570(.A1(new_n639), .A2(new_n657), .A3(new_n725), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n635), .A2(G472), .B1(new_n749), .B2(new_n590), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n746), .A2(new_n757), .A3(new_n687), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  NOR2_X1   g574(.A1(new_n741), .A2(new_n752), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n620), .A2(new_n629), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n442), .A2(new_n447), .A3(new_n444), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n595), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n757), .A4(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n493), .A2(new_n593), .A3(new_n757), .A4(new_n764), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT107), .B(G131), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G33));
  XOR2_X1   g587(.A(new_n695), .B(KEYINPUT108), .Z(new_n774));
  NAND3_X1  g588(.A1(new_n742), .A2(new_n764), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n657), .A2(new_n344), .A3(new_n271), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n636), .A2(new_n637), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n779), .A2(KEYINPUT111), .A3(new_n780), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n687), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n777), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n777), .A3(new_n787), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n626), .A2(new_n628), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT45), .ZN(new_n793));
  OAI21_X1  g607(.A(G469), .B1(new_n792), .B2(KEYINPUT45), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n597), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT109), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n795), .A2(new_n799), .A3(KEYINPUT46), .A4(new_n796), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n731), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  INV_X1    g616(.A(new_n795), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n803), .B2(new_n597), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n797), .A2(KEYINPUT109), .B1(new_n596), .B2(new_n619), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT110), .B1(new_n806), .B2(new_n800), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n594), .B(new_n700), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n763), .ZN(new_n810));
  OAI211_X1 g624(.A(KEYINPUT112), .B(new_n810), .C1(new_n786), .C2(new_n787), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n786), .B2(new_n787), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n791), .A2(new_n809), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  OAI21_X1  g630(.A(new_n594), .B1(new_n805), .B2(new_n807), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT47), .B(new_n594), .C1(new_n805), .C2(new_n807), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n493), .A2(new_n593), .A3(new_n726), .A4(new_n763), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  AOI21_X1  g638(.A(new_n657), .B1(new_n344), .B2(new_n271), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n639), .A2(new_n670), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n446), .A2(new_n334), .A3(new_n448), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n493), .A3(new_n638), .A4(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n689), .B(new_n829), .C1(new_n450), .C2(new_n631), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n747), .A2(new_n755), .A3(new_n734), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(new_n744), .A3(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n630), .A2(new_n488), .A3(new_n686), .A4(new_n725), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n713), .A2(new_n835), .A3(new_n754), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n698), .A2(new_n728), .A3(new_n759), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n728), .A2(new_n698), .A3(new_n759), .A4(new_n836), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n323), .A2(new_n669), .A3(new_n694), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n845), .A2(new_n724), .A3(new_n846), .A4(new_n763), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n593), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n775), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n764), .A2(new_n757), .A3(new_n687), .A4(new_n758), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT116), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n834), .A2(new_n771), .A3(new_n842), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT53), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n832), .B1(new_n740), .B2(new_n743), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n771), .A2(new_n855), .A3(new_n852), .A4(new_n831), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n837), .B2(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n839), .A2(new_n862), .A3(new_n840), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT118), .B1(new_n839), .B2(new_n840), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n839), .A2(new_n862), .A3(new_n840), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n839), .B2(new_n840), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(KEYINPUT54), .B(new_n854), .C1(new_n858), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n856), .A2(new_n857), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n856), .A2(new_n857), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n869), .A3(new_n870), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT54), .A4(new_n854), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n744), .A2(new_n833), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n830), .A2(new_n870), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n771), .A2(new_n852), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(new_n885), .A3(new_n864), .A4(new_n868), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  INV_X1    g701(.A(new_n842), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n870), .B1(new_n856), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n873), .A2(new_n878), .A3(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n732), .A2(new_n763), .A3(new_n328), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n779), .A2(new_n780), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n761), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT48), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n714), .A2(new_n493), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n639), .A3(new_n657), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n781), .A2(new_n328), .A3(new_n752), .A4(new_n751), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n746), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n325), .A2(new_n895), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n639), .A2(new_n657), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n758), .A2(new_n687), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n896), .A2(new_n901), .B1(new_n893), .B2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n898), .A2(new_n448), .A3(new_n708), .A4(new_n733), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT50), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n730), .A2(new_n731), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n595), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n819), .A2(new_n820), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n898), .A2(new_n810), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n909), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n900), .B1(new_n915), .B2(KEYINPUT51), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT51), .B(new_n904), .C1(new_n907), .C2(new_n908), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n912), .B2(KEYINPUT122), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n891), .A2(new_n921), .B1(G952), .B2(G953), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n752), .A2(new_n448), .A3(new_n595), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT114), .Z(new_n924));
  XOR2_X1   g738(.A(new_n910), .B(KEYINPUT49), .Z(new_n925));
  NOR3_X1   g739(.A1(new_n925), .A2(new_n713), .A3(new_n778), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n926), .A3(new_n708), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n194), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n771), .A2(new_n852), .A3(new_n884), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n881), .B2(new_n882), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n932), .A2(new_n869), .B1(new_n870), .B2(new_n853), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n273), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT56), .B1(new_n934), .B2(new_n441), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n420), .A2(new_n421), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n371), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n930), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n935), .B2(new_n938), .ZN(G51));
  NOR3_X1   g754(.A1(new_n933), .A2(new_n273), .A3(new_n795), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n597), .B(KEYINPUT57), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n887), .B1(new_n886), .B2(new_n889), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n614), .ZN(new_n946));
  INV_X1    g760(.A(new_n618), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n941), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT123), .B1(new_n950), .B2(new_n929), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n886), .A2(new_n889), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n890), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n948), .B1(new_n955), .B2(new_n942), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n952), .B(new_n930), .C1(new_n956), .C2(new_n941), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n951), .A2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n268), .A2(new_n246), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n929), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n311), .B1(new_n647), .B2(KEYINPUT99), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n651), .A2(new_n966), .B1(new_n644), .B2(new_n645), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT33), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI221_X1 g783(.A(new_n965), .B1(new_n969), .B2(new_n642), .C1(new_n943), .C2(new_n944), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n930), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n891), .A2(new_n965), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n654), .ZN(G63));
  AND2_X1   g787(.A1(new_n684), .A2(new_n685), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT124), .B1(new_n953), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n979), .B(new_n976), .C1(new_n886), .C2(new_n889), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n974), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n933), .B2(new_n976), .ZN(new_n982));
  INV_X1    g796(.A(new_n484), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n977), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n981), .A2(new_n985), .A3(new_n930), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n981), .A2(new_n985), .A3(KEYINPUT61), .A4(new_n930), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(G66));
  INV_X1    g804(.A(G224), .ZN(new_n991));
  OAI21_X1  g805(.A(G953), .B1(new_n333), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n834), .B2(new_n222), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n936), .B1(G898), .B2(new_n194), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT125), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G69));
  XNOR2_X1  g810(.A(new_n576), .B(new_n239), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(new_n222), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n809), .A2(new_n754), .A3(new_n761), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n823), .A2(new_n771), .A3(new_n775), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n728), .A2(new_n698), .A3(new_n759), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT126), .B1(new_n815), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n814), .A2(new_n789), .A3(new_n811), .A4(new_n790), .ZN(new_n1006));
  OAI211_X1 g820(.A(KEYINPUT126), .B(new_n1004), .C1(new_n1006), .C2(new_n808), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1002), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n999), .B1(new_n1009), .B2(new_n222), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n742), .A2(new_n700), .A3(new_n764), .A4(new_n827), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n716), .A2(new_n1004), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n716), .A2(KEYINPUT62), .A3(new_n1004), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n815), .A2(new_n823), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n997), .B1(new_n1019), .B2(new_n194), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1010), .A2(new_n1012), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n999), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1004), .B1(new_n1006), .B2(new_n808), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1001), .B1(new_n1026), .B2(new_n1007), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1023), .B1(new_n1027), .B2(new_n194), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1011), .B1(new_n1028), .B2(new_n1020), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1022), .A2(new_n1029), .ZN(G72));
  NAND4_X1  g844(.A1(new_n815), .A2(new_n823), .A3(new_n834), .A4(new_n1018), .ZN(new_n1031));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  AND3_X1   g847(.A1(new_n1031), .A2(KEYINPUT127), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(KEYINPUT127), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1035));
  INV_X1    g849(.A(new_n709), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n577), .A2(new_n540), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n1002), .B(new_n834), .C1(new_n1005), .C2(new_n1008), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1038), .B1(new_n1039), .B2(new_n1033), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n876), .A2(new_n854), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1036), .A2(new_n1033), .A3(new_n1038), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n930), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1037), .A2(new_n1040), .A3(new_n1043), .ZN(G57));
endmodule


