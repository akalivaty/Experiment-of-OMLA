//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AND2_X1   g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n215), .B1(new_n202), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n214), .B(new_n217), .C1(G87), .C2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G97), .A2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G77), .A2(G244), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT67), .B(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n201), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n213), .B(new_n227), .C1(new_n235), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G250), .B(G257), .Z(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  AND2_X1   g0055(.A1(KEYINPUT69), .A2(G1), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT69), .A2(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n230), .A2(new_n231), .A3(new_n260), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n259), .A2(new_n202), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT8), .B(G58), .Z(new_n263));
  NAND2_X1  g0063(.A1(new_n234), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n234), .A2(new_n267), .A3(KEYINPUT70), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT70), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G20), .B2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G150), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n203), .A2(KEYINPUT71), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NOR3_X1   g0074(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(new_n234), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n266), .A2(new_n272), .A3(new_n273), .A4(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n262), .B1(new_n277), .B2(new_n261), .ZN(new_n278));
  OAI211_X1 g0078(.A(G13), .B(G20), .C1(new_n256), .C2(new_n257), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n202), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(KEYINPUT73), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT73), .B1(new_n278), .B2(new_n281), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT9), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G222), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G223), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n230), .A2(new_n231), .B1(G33), .B2(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(G77), .C2(new_n288), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT68), .B(G45), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(G274), .C1(new_n296), .C2(G41), .ZN(new_n297));
  INV_X1    g0097(.A(G45), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT69), .A2(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT69), .A2(G1), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(G41), .B1(new_n256), .B2(new_n257), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n294), .B(new_n297), .C1(new_n305), .C2(new_n216), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n277), .A2(new_n261), .ZN(new_n309));
  INV_X1    g0109(.A(new_n262), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n281), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n282), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n306), .A2(G200), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n285), .A2(new_n308), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT10), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n306), .A2(G179), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n306), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n311), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n268), .A2(new_n270), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n202), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT67), .A2(G68), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT67), .A2(G68), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n327), .A2(new_n234), .B1(new_n328), .B2(new_n264), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n261), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT11), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n280), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n279), .A2(G68), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(KEYINPUT12), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NOR4_X1   g0136(.A1(new_n280), .A2(new_n259), .A3(new_n336), .A4(new_n261), .ZN(new_n337));
  OR3_X1    g0137(.A1(new_n332), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI211_X1 g0140(.A(G226), .B(new_n290), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n288), .A2(KEYINPUT74), .A3(G226), .A4(new_n290), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(G232), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n293), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n303), .A2(G238), .A3(new_n304), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n297), .A4(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n343), .B2(new_n344), .ZN(new_n353));
  INV_X1    g0153(.A(new_n293), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n297), .B(new_n351), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT13), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n338), .B1(new_n357), .B2(G200), .ZN(new_n358));
  INV_X1    g0158(.A(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G190), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n318), .A2(new_n322), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT77), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n201), .B1(new_n327), .B2(G58), .ZN(new_n365));
  INV_X1    g0165(.A(G159), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n365), .A2(new_n234), .B1(new_n323), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n286), .A2(new_n234), .A3(new_n287), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n339), .A2(new_n340), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n234), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n223), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n364), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n368), .A2(new_n369), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n371), .B2(new_n234), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G58), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n236), .B1(new_n223), .B2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(G20), .B1(G159), .B2(new_n271), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n380), .A3(KEYINPUT16), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n374), .A2(new_n381), .A3(new_n261), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT8), .B(G58), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n259), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n280), .A2(new_n261), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n263), .A2(new_n258), .A3(KEYINPUT76), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n280), .A2(new_n384), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT69), .B(G1), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G45), .ZN(new_n394));
  INV_X1    g0194(.A(G41), .ZN(new_n395));
  OAI211_X1 g0195(.A(G1), .B(G13), .C1(new_n267), .C2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n394), .A2(G232), .A3(new_n396), .A4(new_n304), .ZN(new_n397));
  NOR2_X1   g0197(.A1(G223), .A2(G1698), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n286), .B2(new_n287), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n216), .A2(G1698), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(G33), .B2(G87), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n397), .B(new_n297), .C1(new_n401), .C2(new_n354), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n293), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(G179), .A3(new_n397), .A4(new_n297), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n392), .A2(KEYINPUT18), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT18), .B1(new_n392), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n363), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n230), .A2(new_n231), .A3(new_n260), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n336), .B1(new_n370), .B2(new_n372), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n367), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n390), .B1(new_n417), .B2(new_n374), .ZN(new_n418));
  INV_X1    g0218(.A(new_n409), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n392), .A2(KEYINPUT18), .A3(new_n409), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(KEYINPUT77), .A3(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n402), .A2(new_n307), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n402), .A2(G200), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n382), .A2(new_n423), .A3(new_n391), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT17), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n412), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n259), .A2(new_n328), .A3(new_n261), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n323), .A2(new_n384), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n431), .A2(new_n264), .B1(new_n234), .B2(new_n328), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n261), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n429), .B1(G77), .B2(new_n279), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n288), .A2(G238), .A3(G1698), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n288), .A2(G232), .A3(new_n290), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n206), .C2(new_n288), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n293), .ZN(new_n440));
  INV_X1    g0240(.A(G244), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n297), .C1(new_n441), .C2(new_n305), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n442), .A2(G179), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n320), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n436), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(G200), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n307), .B2(new_n442), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n436), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT14), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n352), .A2(new_n356), .A3(G179), .ZN(new_n450));
  NAND2_X1  g0250(.A1(KEYINPUT75), .A2(G169), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(new_n450), .C1(new_n359), .C2(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n332), .A2(new_n335), .A3(new_n337), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n352), .B2(new_n356), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(KEYINPUT14), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR4_X1   g0256(.A1(new_n362), .A2(new_n427), .A3(new_n448), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G116), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G20), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n234), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n234), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n461), .A2(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT22), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(new_n286), .B2(new_n287), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(G87), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n234), .B(G87), .C1(new_n339), .C2(new_n340), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(KEYINPUT22), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT88), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT88), .B(new_n466), .C1(new_n469), .C2(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(KEYINPUT24), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n261), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT89), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(KEYINPUT89), .A3(new_n261), .A4(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G33), .B1(new_n256), .B2(new_n257), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n414), .A2(new_n279), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n414), .A2(KEYINPUT78), .A3(new_n279), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n279), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT25), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT5), .B(G41), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n302), .B1(new_n301), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G257), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n498));
  OAI211_X1 g0298(.A(G250), .B(new_n290), .C1(new_n339), .C2(new_n340), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G294), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(G264), .A2(new_n497), .B1(new_n501), .B2(new_n293), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n301), .A2(G274), .A3(new_n496), .A4(new_n396), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(KEYINPUT90), .A3(G179), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT90), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n293), .ZN(new_n506));
  XOR2_X1   g0306(.A(KEYINPUT5), .B(G41), .Z(new_n507));
  OAI211_X1 g0307(.A(G264), .B(new_n396), .C1(new_n394), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n509), .B2(G169), .ZN(new_n510));
  INV_X1    g0310(.A(G179), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n504), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT91), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT91), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n515), .B(new_n504), .C1(new_n510), .C2(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n495), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n489), .A2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n521), .A2(new_n205), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n234), .B1(new_n328), .B2(new_n323), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n206), .B1(new_n370), .B2(new_n372), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n261), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n520), .B(new_n527), .C1(G97), .C2(new_n279), .ZN(new_n528));
  OAI211_X1 g0328(.A(G244), .B(new_n290), .C1(new_n339), .C2(new_n340), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n293), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n497), .A2(G257), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n503), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n320), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n535), .A2(new_n293), .B1(G257), .B2(new_n497), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n511), .A3(new_n503), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n528), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n489), .A2(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT82), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n489), .A2(new_n545), .A3(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n224), .A2(new_n290), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n441), .A2(G1698), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n339), .C2(new_n340), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n460), .ZN(new_n551));
  AOI22_X1  g0351(.A1(G250), .A2(new_n303), .B1(new_n551), .B2(new_n293), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT80), .ZN(new_n553));
  OAI211_X1 g0353(.A(G45), .B(G274), .C1(new_n256), .C2(new_n257), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n302), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n301), .A2(KEYINPUT80), .A3(G274), .A4(new_n396), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G190), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n468), .A2(G68), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n234), .B1(new_n347), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G87), .B2(new_n207), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n264), .B2(new_n205), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n261), .B1(new_n280), .B2(new_n431), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n547), .A2(new_n560), .A3(new_n561), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT79), .B1(new_n538), .B2(new_n307), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n523), .A2(new_n521), .ZN(new_n571));
  INV_X1    g0371(.A(new_n522), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n271), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n375), .B2(new_n376), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n414), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n205), .B1(new_n487), .B2(new_n488), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n279), .A2(G97), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n538), .A2(G200), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT79), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n540), .A2(new_n581), .A3(G190), .A4(new_n503), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n570), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n552), .A2(G179), .A3(new_n557), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n320), .B1(new_n552), .B2(new_n557), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT81), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n558), .A2(G169), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n552), .A2(G179), .A3(new_n557), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n431), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n489), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n568), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n586), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n542), .A2(new_n569), .A3(new_n583), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n509), .A2(G190), .ZN(new_n596));
  INV_X1    g0396(.A(G200), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n509), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n483), .A2(new_n494), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n386), .A2(G116), .A3(new_n484), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n279), .A2(KEYINPUT84), .A3(G116), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT84), .B1(new_n279), .B2(G116), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G20), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n533), .B(new_n234), .C1(G33), .C2(new_n205), .ZN(new_n607));
  OR2_X1    g0407(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n261), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n601), .B(new_n604), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(G264), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n614));
  OAI211_X1 g0414(.A(G257), .B(new_n290), .C1(new_n339), .C2(new_n340), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n286), .A2(G303), .A3(new_n287), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT83), .A4(new_n616), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n293), .A3(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n554), .A2(new_n507), .A3(new_n302), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(G270), .B2(new_n497), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n613), .A2(new_n624), .A3(G169), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT86), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT86), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n613), .A2(new_n624), .A3(new_n628), .A4(G169), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n627), .B(new_n320), .C1(new_n621), .C2(new_n623), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n624), .A2(new_n511), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n613), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(G200), .ZN(new_n634));
  INV_X1    g0434(.A(new_n613), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n634), .B(new_n635), .C1(new_n307), .C2(new_n624), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n630), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n519), .A2(new_n595), .A3(new_n600), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n458), .A2(new_n638), .ZN(G372));
  AOI21_X1  g0439(.A(new_n493), .B1(new_n481), .B2(new_n482), .ZN(new_n640));
  INV_X1    g0440(.A(new_n513), .ZN(new_n641));
  OR3_X1    g0441(.A1(new_n640), .A2(KEYINPUT93), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n630), .A2(new_n633), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT93), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n545), .B1(new_n489), .B2(G87), .ZN(new_n647));
  INV_X1    g0447(.A(G87), .ZN(new_n648));
  AOI211_X1 g0448(.A(KEYINPUT82), .B(new_n648), .C1(new_n487), .C2(new_n488), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n561), .B(new_n568), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT92), .B1(new_n584), .B2(new_n585), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT92), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n587), .A2(new_n653), .A3(new_n589), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n651), .A2(new_n560), .B1(new_n655), .B2(new_n593), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n583), .A2(new_n542), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n600), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n593), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n528), .A2(new_n539), .A3(new_n541), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n569), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(new_n661), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n569), .A2(new_n662), .A3(new_n594), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(KEYINPUT26), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n660), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n457), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT94), .ZN(new_n670));
  INV_X1    g0470(.A(new_n322), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n420), .A2(new_n421), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT95), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n445), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n436), .A2(new_n443), .A3(KEYINPUT95), .A4(new_n444), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n456), .B1(new_n676), .B2(new_n361), .ZN(new_n677));
  INV_X1    g0477(.A(new_n426), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n671), .B1(new_n679), .B2(new_n318), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n670), .A2(new_n680), .ZN(G369));
  NOR2_X1   g0481(.A1(new_n640), .A2(new_n517), .ZN(new_n682));
  AOI211_X1 g0482(.A(new_n493), .B(new_n598), .C1(new_n481), .C2(new_n482), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G13), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G20), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n393), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n684), .B1(new_n640), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n519), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n643), .A2(new_n693), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n613), .A2(new_n692), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n637), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n644), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n692), .B1(new_n642), .B2(new_n645), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n684), .B2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n211), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n237), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n665), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n643), .B1(new_n495), .B2(new_n518), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n658), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n693), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n720), .B(new_n661), .C1(KEYINPUT26), .C2(new_n663), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n646), .B2(new_n659), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n692), .ZN(new_n723));
  XNOR2_X1  g0523(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n684), .A2(new_n595), .A3(new_n637), .A4(new_n693), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n540), .A2(new_n552), .A3(new_n557), .ZN(new_n728));
  INV_X1    g0528(.A(new_n509), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n728), .A2(new_n632), .A3(KEYINPUT30), .A4(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(G179), .A3(new_n623), .A4(new_n621), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n559), .A2(new_n540), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n540), .A2(new_n503), .B1(new_n623), .B2(new_n621), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n511), .A3(new_n558), .A4(new_n509), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n730), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n692), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n740), .A3(new_n692), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n726), .B1(new_n727), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n725), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n714), .B1(new_n746), .B2(G1), .ZN(G364));
  NAND2_X1  g0547(.A1(new_n686), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n710), .A2(G1), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n703), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n701), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n233), .B1(G20), .B2(new_n320), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n708), .A2(new_n371), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G355), .A2(new_n759), .B1(new_n605), .B2(new_n708), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n371), .A2(new_n211), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT98), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n763), .B1(new_n238), .B2(new_n296), .C1(new_n298), .C2(new_n254), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n758), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n234), .A2(new_n511), .A3(KEYINPUT99), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT99), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G20), .B2(G179), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n307), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT100), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n769), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n307), .A2(new_n597), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n775), .A2(G322), .B1(G326), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n597), .A2(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(G311), .ZN(new_n786));
  INV_X1    g0586(.A(G303), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n234), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n777), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(new_n307), .A3(new_n597), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n288), .B1(new_n792), .B2(G329), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n307), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n234), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n788), .A2(new_n781), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n780), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n796), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n775), .A2(G58), .B1(G97), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n785), .A2(G77), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n791), .A2(new_n366), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n806), .A2(KEYINPUT32), .B1(new_n336), .B2(new_n782), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n800), .A2(new_n206), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(KEYINPUT32), .ZN(new_n810));
  INV_X1    g0610(.A(new_n789), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G87), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n779), .A2(G50), .ZN(new_n813));
  AND4_X1   g0613(.A1(new_n288), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n803), .A2(new_n804), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n749), .B(new_n765), .C1(new_n816), .C2(new_n753), .ZN(new_n817));
  INV_X1    g0617(.A(new_n756), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n701), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n752), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  AOI22_X1  g0621(.A1(new_n775), .A2(G143), .B1(G159), .B2(new_n785), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  INV_X1    g0623(.A(G150), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n778), .B1(new_n782), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT103), .Z(new_n826));
  NAND2_X1  g0626(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT34), .Z(new_n828));
  OAI22_X1  g0628(.A1(new_n789), .A2(new_n202), .B1(new_n800), .B2(new_n336), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n828), .A2(new_n371), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n378), .B2(new_n796), .C1(new_n831), .C2(new_n791), .ZN(new_n832));
  INV_X1    g0632(.A(G311), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n791), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n774), .A2(new_n794), .B1(new_n787), .B2(new_n778), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G116), .B2(new_n785), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n800), .A2(new_n648), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G97), .B2(new_n802), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT102), .B(G283), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n371), .B1(new_n782), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G107), .B2(new_n811), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n836), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n832), .B1(new_n834), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n753), .A2(new_n754), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n844), .A2(new_n753), .B1(new_n328), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n750), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT104), .Z(new_n848));
  NAND4_X1  g0648(.A1(new_n674), .A2(new_n436), .A3(new_n675), .A4(new_n692), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n436), .A2(new_n692), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n448), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n848), .B1(new_n755), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n723), .B(new_n853), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n744), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT106), .Z(new_n857));
  OR2_X1    g0657(.A1(new_n855), .A2(new_n744), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n750), .B1(new_n858), .B2(KEYINPUT105), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(KEYINPUT105), .C2(new_n858), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(G384));
  OAI211_X1 g0661(.A(new_n235), .B(G116), .C1(new_n573), .C2(KEYINPUT35), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT107), .Z(new_n863));
  INV_X1    g0663(.A(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n864), .B2(new_n524), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT36), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n328), .B(new_n237), .C1(new_n327), .C2(G58), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n336), .A2(G50), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n685), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n358), .A2(new_n360), .B1(new_n338), .B2(new_n692), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT108), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT108), .B1(new_n452), .B2(new_n455), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n456), .A2(new_n692), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n668), .A2(new_n693), .A3(new_n853), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n445), .A2(new_n692), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n381), .A2(new_n261), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n391), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n690), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n427), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n392), .B1(new_n409), .B2(new_n883), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n425), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n882), .A2(new_n409), .ZN(new_n890));
  INV_X1    g0690(.A(new_n425), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n892), .B2(new_n888), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n879), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n420), .A2(new_n421), .A3(new_n690), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n423), .A4(new_n424), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT17), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n425), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n902), .B(new_n904), .C1(new_n410), .C2(new_n411), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n418), .A2(new_n690), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n419), .A2(new_n690), .B1(new_n382), .B2(new_n391), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n907), .B2(new_n891), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n905), .A2(new_n906), .B1(new_n908), .B2(new_n889), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT109), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT109), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n908), .A2(new_n889), .ZN(new_n912));
  INV_X1    g0712(.A(new_n906), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n426), .B2(new_n672), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n911), .B(new_n895), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n897), .A2(new_n910), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n901), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n871), .A2(new_n872), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n693), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n899), .A2(new_n900), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n457), .B(new_n719), .C1(new_n723), .C2(new_n724), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n680), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n897), .A2(new_n910), .A3(new_n915), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n742), .B1(new_n638), .B2(new_n692), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n873), .A2(new_n874), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n853), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT40), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n852), .B1(new_n727), .B2(new_n742), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n898), .A2(new_n932), .A3(new_n929), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n457), .A3(new_n928), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(G330), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n457), .A2(new_n743), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n936), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n926), .A2(new_n941), .B1(new_n393), .B2(new_n686), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT110), .Z(new_n943));
  AND2_X1   g0743(.A1(new_n926), .A2(new_n941), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n866), .B1(new_n393), .B2(new_n869), .C1(new_n943), .C2(new_n944), .ZN(G367));
  NAND2_X1  g0745(.A1(new_n775), .A2(G303), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n789), .A2(new_n605), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n947), .A2(KEYINPUT46), .B1(new_n792), .B2(G317), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n785), .A2(new_n839), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n946), .A2(new_n371), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n947), .A2(KEYINPUT46), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n778), .A2(new_n833), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n796), .A2(new_n206), .ZN(new_n953));
  NOR4_X1   g0753(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n205), .B2(new_n800), .C1(new_n794), .C2(new_n782), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT112), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n371), .B1(new_n775), .B2(G150), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n779), .A2(G143), .ZN(new_n958));
  INV_X1    g0758(.A(new_n785), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n202), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n782), .A2(new_n366), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n800), .A2(new_n328), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n823), .A2(new_n791), .B1(new_n789), .B2(new_n378), .ZN(new_n963));
  NOR4_X1   g0763(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n796), .A2(new_n336), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n957), .A2(new_n958), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n956), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n753), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n547), .A2(new_n568), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n692), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n656), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n661), .B2(new_n972), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(new_n818), .ZN(new_n975));
  INV_X1    g0775(.A(new_n763), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n757), .B1(new_n211), .B2(new_n431), .C1(new_n976), .C2(new_n247), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n970), .A2(new_n750), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n684), .A2(new_n697), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n657), .B1(new_n579), .B2(new_n693), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT42), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n542), .B1(new_n982), .B2(new_n519), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n985), .A2(new_n693), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n980), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT111), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(new_n989), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n662), .A2(new_n692), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n982), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n704), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n992), .B(new_n996), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n706), .A2(new_n994), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT45), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n706), .A2(new_n994), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n704), .A3(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n698), .A2(new_n703), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n1003), .A2(new_n704), .A3(new_n981), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n745), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(G1), .B(new_n748), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n979), .B1(new_n997), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(G387));
  NAND2_X1  g0810(.A1(new_n748), .A2(G1), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n296), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n763), .B1(new_n244), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n759), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n711), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT50), .B1(new_n384), .B2(G50), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n711), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n384), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1018), .A2(G45), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n336), .B2(new_n328), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n708), .A2(new_n206), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n758), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n775), .A2(G50), .B1(G68), .B2(new_n785), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n288), .B1(new_n205), .B2(new_n800), .C1(new_n778), .C2(new_n366), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n796), .A2(new_n431), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n791), .A2(new_n824), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n789), .A2(new_n328), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1025), .B(new_n1030), .C1(new_n384), .C2(new_n782), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n779), .A2(G322), .B1(new_n785), .B2(G303), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n833), .B2(new_n782), .C1(new_n774), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT48), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n794), .B2(new_n789), .C1(new_n796), .C2(new_n840), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT49), .Z(new_n1037));
  AOI21_X1  g0837(.A(new_n288), .B1(new_n792), .B2(G326), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n605), .B2(new_n800), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1031), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1024), .B1(new_n1040), .B2(new_n753), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n750), .C1(new_n695), .C2(new_n818), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1004), .A2(new_n746), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n709), .B1(new_n1004), .B2(new_n746), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1012), .B(new_n1042), .C1(new_n1043), .C2(new_n1044), .ZN(G393));
  OAI221_X1 g0845(.A(new_n757), .B1(new_n205), .B2(new_n211), .C1(new_n976), .C2(new_n251), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n750), .B(new_n1046), .C1(new_n994), .C2(new_n818), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n774), .A2(new_n366), .B1(new_n824), .B2(new_n778), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT51), .Z(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G77), .B2(new_n802), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n792), .A2(G143), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n371), .B1(new_n783), .B2(G50), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n789), .A2(new_n223), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n837), .B(new_n1053), .C1(new_n785), .C2(new_n263), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n774), .A2(new_n833), .B1(new_n1033), .B2(new_n778), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  AOI211_X1 g0857(.A(new_n288), .B(new_n1057), .C1(G322), .C2(new_n792), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n782), .A2(new_n787), .B1(new_n605), .B2(new_n796), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n808), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n794), .C2(new_n959), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n840), .A2(new_n789), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1047), .B1(new_n1063), .B2(new_n753), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1002), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n704), .B1(new_n999), .B2(new_n1001), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n1067), .B2(new_n1011), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1043), .A2(new_n1002), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1067), .B2(new_n1043), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1070), .B2(new_n710), .ZN(G390));
  NAND3_X1  g0871(.A1(new_n743), .A2(new_n853), .A3(new_n929), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT113), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n718), .A2(new_n693), .A3(new_n853), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n878), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n929), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n897), .A2(new_n910), .A3(new_n915), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n920), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1074), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n875), .B1(new_n1075), .B2(new_n878), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n920), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1081), .A2(new_n1082), .A3(KEYINPUT113), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n722), .A2(new_n692), .A3(new_n852), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n929), .B1(new_n1085), .B2(new_n877), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n918), .B1(new_n1086), .B2(new_n920), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1073), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n901), .A2(new_n917), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n879), .B2(new_n921), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1077), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT113), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1093), .A3(new_n1072), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n924), .A2(new_n680), .A3(new_n939), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n876), .A2(new_n878), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n929), .B1(new_n743), .B2(new_n853), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT114), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1072), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n928), .A2(G330), .A3(new_n853), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1101), .A2(new_n1099), .A3(new_n875), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1097), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n875), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n743), .B(new_n853), .C1(KEYINPUT115), .C2(new_n929), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n878), .A4(new_n1075), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1096), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1095), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1088), .A2(new_n1108), .A3(new_n1094), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n709), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n754), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n783), .A2(G137), .B1(G159), .B2(new_n802), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n800), .A2(new_n202), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n371), .B(new_n1115), .C1(G125), .C2(new_n792), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1114), .B(new_n1116), .C1(new_n1117), .C2(new_n778), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  NAND2_X1  g0919(.A1(new_n785), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n811), .A2(G150), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1120), .B1(KEYINPUT53), .B2(new_n1121), .C1(new_n774), .C2(new_n831), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1118), .B(new_n1122), .C1(KEYINPUT53), .C2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n774), .A2(new_n605), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n288), .B1(new_n785), .B2(G97), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n328), .B2(new_n796), .C1(new_n206), .C2(new_n782), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n778), .A2(new_n799), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n812), .B1(new_n800), .B2(new_n336), .C1(new_n794), .C2(new_n791), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n753), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n845), .A2(new_n384), .ZN(new_n1131));
  AND4_X1   g0931(.A1(new_n750), .A2(new_n1113), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1095), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n1011), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1112), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1112), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(new_n1096), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1111), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n322), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n283), .A2(new_n284), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n883), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n318), .A2(new_n322), .A3(new_n1147), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1078), .A2(new_n933), .A3(new_n929), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n930), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT40), .B1(new_n896), .B2(new_n897), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1155), .A2(KEYINPUT40), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1154), .B1(new_n1158), .B2(new_n726), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1154), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n935), .A2(G330), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n923), .A2(new_n1142), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1160), .B1(new_n935), .B2(G330), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n726), .B(new_n1154), .C1(new_n931), .C2(new_n934), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT120), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n923), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1159), .A2(new_n1142), .A3(new_n1161), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1141), .A2(KEYINPUT57), .A3(new_n1162), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n709), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT121), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT119), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(new_n923), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1141), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1169), .A2(KEYINPUT121), .A3(new_n709), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1172), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1174), .A2(new_n1011), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n774), .A2(new_n206), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT117), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n800), .A2(new_n378), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1029), .B(new_n1183), .C1(new_n785), .C2(new_n591), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n395), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G283), .B2(new_n792), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n288), .B(new_n965), .C1(new_n783), .C2(G97), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n605), .C2(new_n778), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT58), .Z(new_n1189));
  OAI21_X1  g0989(.A(new_n202), .B1(new_n339), .B2(G41), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G125), .A2(new_n779), .B1(new_n783), .B2(G132), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G137), .B2(new_n785), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n802), .A2(G150), .B1(new_n811), .B2(new_n1119), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n1117), .C2(new_n774), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G33), .B1(new_n1195), .B2(KEYINPUT59), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT118), .B(G124), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G41), .B1(new_n792), .B2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(new_n366), .C2(new_n800), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1190), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n753), .B1(new_n1189), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n845), .A2(new_n202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n749), .B1(new_n1154), .B2(new_n754), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1180), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1179), .A2(new_n1207), .ZN(G375));
  NAND3_X1  g1008(.A1(new_n1103), .A2(new_n1096), .A3(new_n1107), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1109), .A2(new_n1006), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n875), .A2(new_n754), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n778), .A2(new_n794), .B1(new_n787), .B2(new_n791), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n959), .A2(new_n206), .B1(new_n782), .B2(new_n605), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n288), .B(new_n1212), .C1(new_n1213), .C2(KEYINPUT123), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(KEYINPUT123), .B2(new_n1213), .C1(new_n799), .C2(new_n774), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n789), .A2(new_n205), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(new_n962), .A3(new_n1027), .A4(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n775), .A2(G137), .B1(G50), .B2(new_n802), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n783), .A2(new_n1119), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n378), .C2(new_n800), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n791), .A2(new_n1117), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n959), .A2(new_n824), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n288), .B1(new_n366), .B2(new_n789), .C1(new_n778), .C2(new_n831), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n753), .B1(new_n1217), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n845), .A2(new_n336), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n750), .A2(new_n1211), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1011), .B(KEYINPUT122), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1210), .A2(new_n1230), .ZN(G381));
  NOR2_X1   g1031(.A1(G375), .A2(new_n1135), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1233), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1234), .B2(new_n1237), .ZN(G407));
  OAI211_X1 g1039(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  NAND3_X1  g1040(.A1(new_n1179), .A2(G378), .A3(new_n1207), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1168), .A2(new_n1162), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1229), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1205), .C1(new_n1175), .C2(new_n1007), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1135), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1209), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1209), .A2(new_n1251), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n709), .A3(new_n1109), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G384), .A2(new_n1230), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1230), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n854), .A3(new_n860), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1247), .A2(new_n1250), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1249), .A2(G2897), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1258), .B(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1246), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1176), .B1(new_n1111), .B2(new_n1140), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1171), .B(new_n710), .C1(new_n1242), .C2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT121), .B1(new_n1169), .B2(new_n709), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1206), .B1(new_n1269), .B2(new_n1177), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1265), .B1(new_n1270), .B2(G378), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1264), .B1(new_n1271), .B2(new_n1249), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1247), .A2(new_n1273), .A3(new_n1259), .A4(new_n1250), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1261), .A2(new_n1262), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n820), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1009), .A2(G390), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1009), .A2(G390), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT126), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n1276), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  OR3_X1    g1084(.A1(new_n1009), .A2(KEYINPUT127), .A3(G390), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1276), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT127), .B1(new_n1009), .B2(G390), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1285), .A2(new_n1277), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1275), .A2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT125), .B1(new_n1271), .B2(new_n1249), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1247), .A2(new_n1292), .A3(new_n1250), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1264), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1260), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1259), .A4(new_n1250), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1294), .A2(new_n1295), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1290), .A2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1245), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1241), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1259), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1241), .A3(new_n1258), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1289), .B(new_n1305), .ZN(G402));
endmodule


