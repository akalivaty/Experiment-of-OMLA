//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT64), .B1(new_n200), .B2(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n198), .A3(G146), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n199), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n204), .A2(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n197), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n202), .B1(new_n198), .B2(G146), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n200), .A2(KEYINPUT64), .A3(G143), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n206), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n208), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n188), .A2(G137), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n190), .A2(G134), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n196), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G116), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n234), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n212), .A2(new_n227), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n196), .A2(new_n225), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n218), .B2(new_n221), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n246), .A2(new_n247), .B1(new_n197), .B2(new_n211), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n204), .A2(new_n215), .B1(new_n220), .B2(new_n208), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT65), .B1(new_n249), .B2(new_n245), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(KEYINPUT67), .A3(new_n239), .A4(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n222), .A2(new_n226), .A3(new_n247), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n250), .A2(new_n252), .A3(new_n239), .A4(new_n212), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n238), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n244), .B1(new_n259), .B2(KEYINPUT28), .ZN(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G237), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT69), .B(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n260), .A2(KEYINPUT71), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n242), .B(KEYINPUT70), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n251), .A2(new_n255), .B1(new_n257), .B2(new_n238), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n275), .B(new_n273), .C1(new_n276), .C2(new_n241), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n251), .A2(KEYINPUT28), .A3(new_n255), .ZN(new_n282));
  INV_X1    g096(.A(new_n271), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n197), .A2(new_n211), .B1(new_n222), .B2(new_n226), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n239), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n241), .B2(new_n240), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n272), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n238), .B1(new_n284), .B2(KEYINPUT30), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT30), .A4(new_n212), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n291), .A2(KEYINPUT66), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(KEYINPUT66), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n283), .B1(new_n294), .B2(new_n256), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n281), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G472), .B1(new_n280), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n253), .A2(new_n254), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n253), .A2(new_n254), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n283), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n248), .A2(new_n303), .A3(KEYINPUT30), .A4(new_n250), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n291), .A2(KEYINPUT66), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n289), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n299), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n271), .B1(new_n251), .B2(new_n255), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n283), .B1(new_n282), .B2(new_n286), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G472), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n298), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n307), .B2(new_n309), .ZN(new_n316));
  NOR4_X1   g130(.A1(new_n316), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n297), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(G234), .B2(new_n281), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT73), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT73), .A3(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n327), .A2(KEYINPUT16), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n200), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n338), .A2(G146), .A3(new_n333), .A4(new_n332), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(KEYINPUT75), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n341), .B(new_n200), .C1(new_n334), .C2(new_n335), .ZN(new_n342));
  INV_X1    g156(.A(G128), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(new_n343), .B2(G119), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT72), .B1(new_n228), .B2(G128), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G110), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(G119), .B(G128), .Z(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT24), .B(G110), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n340), .A2(new_n342), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n200), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n346), .A2(new_n347), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n349), .A2(new_n350), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n339), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT77), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n353), .A2(new_n358), .A3(new_n364), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n281), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n323), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n369), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n366), .A2(new_n281), .A3(new_n367), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n321), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n320), .A2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n366), .B2(new_n367), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n366), .A2(new_n376), .A3(new_n367), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n318), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n218), .A2(new_n221), .A3(new_n324), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n211), .B2(new_n324), .ZN(new_n385));
  INV_X1    g199(.A(G224), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G953), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n385), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G122), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n392));
  OR2_X1    g206(.A1(KEYINPUT81), .A2(G107), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT81), .A2(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n401), .A2(new_n402), .B1(new_n236), .B2(new_n237), .ZN(new_n403));
  AND2_X1   g217(.A1(KEYINPUT81), .A2(G107), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT81), .A2(G107), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n399), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G107), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(new_n392), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n400), .A3(new_n390), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(KEYINPUT4), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n413));
  INV_X1    g227(.A(G113), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n230), .A2(G119), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n413), .A2(new_n417), .B1(new_n233), .B2(new_n235), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n390), .B1(G104), .B2(G107), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n393), .A2(new_n394), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(G104), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n410), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n389), .B1(new_n412), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT85), .B(KEYINPUT6), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n412), .A2(new_n389), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT6), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(new_n424), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n403), .A2(new_n411), .B1(new_n418), .B2(new_n422), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(new_n389), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n412), .A2(new_n423), .ZN(new_n434));
  INV_X1    g248(.A(new_n389), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT84), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n388), .B(new_n426), .C1(new_n430), .C2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n211), .A2(new_n324), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n249), .A2(new_n440), .A3(new_n324), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n384), .A2(KEYINPUT88), .ZN(new_n442));
  INV_X1    g256(.A(new_n387), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n439), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(new_n427), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n449));
  OAI21_X1  g263(.A(G113), .B1(new_n229), .B2(KEYINPUT5), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n413), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n422), .A2(new_n236), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n455));
  INV_X1    g269(.A(new_n418), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n410), .A2(new_n421), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n454), .A2(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n422), .A2(KEYINPUT87), .A3(new_n453), .A4(new_n236), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n389), .B(KEYINPUT8), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n448), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G210), .B1(G237), .B2(G902), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n438), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n438), .B2(new_n463), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n383), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT89), .B(new_n383), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(G110), .B(G140), .Z(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT80), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n266), .A2(G227), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n343), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n204), .A2(new_n478), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n214), .B(new_n199), .C1(new_n201), .C2(new_n203), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n410), .B(new_n421), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n401), .A2(new_n402), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n411), .A2(new_n211), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n197), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n422), .A2(KEYINPUT10), .A3(new_n222), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n457), .A2(new_n249), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n486), .B1(new_n481), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n495), .B(new_n486), .C1(new_n481), .C2(new_n493), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n477), .B(new_n488), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n197), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n477), .B1(new_n501), .B2(new_n488), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n502), .B2(KEYINPUT83), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n481), .A2(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n197), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n491), .B1(new_n505), .B2(new_n495), .ZN(new_n506));
  INV_X1    g320(.A(new_n498), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n477), .A4(new_n488), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G469), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n281), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n514));
  INV_X1    g328(.A(new_n477), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n501), .A2(new_n477), .A3(new_n488), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(G469), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(G469), .A2(G902), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n473), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n469), .A2(new_n470), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n198), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n265), .A2(new_n266), .A3(G143), .A4(G214), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT18), .A3(G131), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n355), .B1(new_n330), .B2(new_n200), .ZN(new_n528));
  NAND2_X1  g342(.A1(KEYINPUT18), .A2(G131), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n195), .B1(new_n524), .B2(new_n525), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n524), .A2(new_n195), .A3(new_n525), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n533), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n536), .A2(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n340), .A2(new_n342), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n532), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G113), .B(G122), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n391), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT90), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n545), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n354), .A2(KEYINPUT19), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n330), .B2(KEYINPUT19), .ZN(new_n550));
  OAI221_X1 g364(.A(new_n339), .B1(G146), .B2(new_n550), .C1(new_n538), .C2(new_n533), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n548), .B1(new_n552), .B2(new_n532), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G475), .A2(G902), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT20), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  XNOR2_X1  g376(.A(G116), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT94), .ZN(new_n564));
  INV_X1    g378(.A(new_n420), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XOR2_X1   g381(.A(G128), .B(G143), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G134), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n230), .A2(KEYINPUT14), .A3(G122), .ZN(new_n570));
  INV_X1    g384(.A(new_n563), .ZN(new_n571));
  OAI211_X1 g385(.A(G107), .B(new_n570), .C1(new_n571), .C2(KEYINPUT14), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT96), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n566), .A2(new_n575), .A3(new_n572), .A4(new_n569), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n198), .A2(G128), .B1(KEYINPUT95), .B2(KEYINPUT13), .ZN(new_n578));
  AND2_X1   g392(.A1(KEYINPUT95), .A2(KEYINPUT13), .ZN(new_n579));
  OAI21_X1  g393(.A(G134), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n568), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n564), .A2(new_n565), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n567), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n471), .A2(new_n319), .A3(G953), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n583), .A3(new_n585), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n562), .B1(new_n589), .B2(new_n281), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n577), .A2(new_n583), .A3(new_n585), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n585), .B1(new_n577), .B2(new_n583), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n281), .B(new_n562), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G953), .ZN(new_n596));
  INV_X1    g410(.A(G952), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(G234), .B2(G237), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n281), .B(new_n266), .C1(G234), .C2(G237), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT21), .B(G898), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n548), .B1(new_n543), .B2(KEYINPUT92), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n607), .B(new_n532), .C1(new_n541), .C2(new_n542), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n547), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT93), .A3(new_n281), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G475), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT93), .B1(new_n609), .B2(new_n281), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n560), .B(new_n605), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n382), .A2(new_n522), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n390), .ZN(G3));
  OAI21_X1  g429(.A(new_n560), .B1(new_n611), .B2(new_n612), .ZN(new_n616));
  AOI21_X1  g430(.A(G478), .B1(new_n589), .B2(new_n281), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n589), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n561), .A2(G902), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n467), .A2(new_n604), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n616), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n316), .B2(G902), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n302), .A2(new_n306), .A3(new_n299), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT31), .B1(new_n294), .B2(new_n308), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n312), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n314), .A3(new_n281), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n627), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n281), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(KEYINPUT98), .A3(G472), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n381), .A3(new_n521), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(new_n391), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  OAI211_X1 g455(.A(new_n560), .B(new_n595), .C1(new_n611), .C2(new_n612), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n604), .A3(new_n467), .ZN(new_n643));
  INV_X1    g457(.A(new_n637), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n396), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n522), .A2(new_n613), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n368), .A2(new_n369), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n372), .A3(new_n322), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n320), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n365), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n359), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n374), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n601), .B1(new_n602), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n631), .A2(KEYINPUT32), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n313), .A2(new_n298), .A3(new_n314), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n288), .A2(new_n295), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n274), .A3(new_n281), .A4(new_n279), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n666), .A2(new_n667), .B1(new_n669), .B2(G472), .ZN(new_n670));
  INV_X1    g484(.A(new_n383), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n438), .A2(new_n463), .ZN(new_n672));
  INV_X1    g486(.A(new_n464), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n438), .A2(new_n463), .A3(new_n464), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n521), .B(new_n676), .C1(new_n373), .C2(new_n655), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n665), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI211_X1 g494(.A(G469), .B(G902), .C1(new_n503), .C2(new_n510), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n518), .A2(new_n519), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n472), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n467), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n318), .A2(new_n657), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n609), .A2(new_n281), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT93), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(G475), .A3(new_n610), .ZN(new_n689));
  INV_X1    g503(.A(new_n664), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n560), .A3(new_n595), .A4(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT102), .B1(new_n685), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n680), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  NOR2_X1   g508(.A1(new_n465), .A2(new_n466), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  INV_X1    g510(.A(new_n595), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n696), .A2(new_n697), .A3(new_n671), .A4(new_n657), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n664), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n521), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n302), .A2(new_n306), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n271), .B2(new_n259), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n704), .B2(G902), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n315), .B2(new_n317), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n698), .A2(new_n616), .A3(new_n702), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NAND3_X1  g522(.A1(new_n616), .A2(new_n624), .A3(new_n690), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n685), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n200), .ZN(G48));
  NAND2_X1  g525(.A1(new_n511), .A2(new_n281), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n472), .A3(new_n513), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n318), .A2(new_n381), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n626), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  INV_X1    g532(.A(new_n379), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n377), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n652), .B1(new_n375), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n713), .A2(new_n472), .A3(new_n513), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n670), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n643), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT104), .B(G116), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G18));
  INV_X1    g540(.A(new_n613), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n467), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n318), .A3(new_n657), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  OAI21_X1  g544(.A(new_n310), .B1(new_n283), .B2(new_n260), .ZN(new_n731));
  NOR2_X1   g545(.A1(G472), .A2(G902), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n627), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n721), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n467), .A2(new_n697), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n722), .A2(new_n604), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n735), .A2(new_n616), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  AOI21_X1  g553(.A(new_n655), .B1(new_n320), .B2(new_n651), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n734), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n728), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n709), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n324), .ZN(G27));
  NAND3_X1  g558(.A1(new_n674), .A2(new_n383), .A3(new_n675), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n683), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n318), .A2(new_n381), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n623), .B1(new_n689), .B2(new_n560), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n748), .A4(new_n690), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n318), .A2(new_n381), .A3(new_n746), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n709), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND2_X1  g568(.A1(new_n747), .A2(new_n665), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(new_n517), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n515), .B2(new_n514), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n519), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT105), .A3(new_n513), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n761), .A2(new_n519), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(KEYINPUT46), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT105), .B1(new_n762), .B2(new_n513), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n473), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n745), .B(KEYINPUT107), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n699), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n636), .A2(new_n740), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT106), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n616), .B2(new_n623), .ZN(new_n774));
  INV_X1    g588(.A(new_n616), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT43), .A3(new_n624), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n772), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n770), .B1(KEYINPUT44), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(KEYINPUT44), .B2(new_n777), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n767), .B2(new_n473), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT47), .B(new_n472), .C1(new_n765), .C2(new_n766), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n745), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n616), .A2(new_n624), .A3(new_n690), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n670), .A3(new_n721), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND3_X1  g603(.A1(new_n624), .A2(new_n383), .A3(new_n472), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n713), .A2(new_n513), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT49), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(KEYINPUT49), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n706), .A2(new_n721), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n775), .A3(new_n696), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n713), .A2(new_n473), .A3(new_n513), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n782), .A2(new_n783), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(new_n769), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n776), .A2(new_n774), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(KEYINPUT112), .A3(new_n601), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT112), .B1(new_n800), .B2(new_n601), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n735), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n799), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n722), .A2(new_n745), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n741), .B(new_n808), .C1(new_n802), .C2(new_n803), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n795), .A2(new_n601), .A3(new_n808), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n775), .A3(new_n623), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n798), .A2(new_n769), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT113), .B1(new_n813), .B2(new_n804), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n807), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n696), .A2(new_n671), .A3(new_n714), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT114), .Z(new_n817));
  OAI211_X1 g631(.A(new_n735), .B(new_n817), .C1(new_n802), .C2(new_n803), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT50), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n600), .B1(new_n810), .B2(new_n748), .ZN(new_n822));
  INV_X1    g636(.A(new_n728), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n804), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n670), .A2(new_n721), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n808), .C1(new_n802), .C2(new_n803), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT48), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(KEYINPUT48), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n812), .B(KEYINPUT51), .C1(new_n804), .C2(new_n813), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n819), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n821), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n807), .A2(new_n812), .A3(new_n814), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n819), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n830), .A2(new_n819), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n829), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT109), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT108), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n595), .A2(new_n664), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n689), .A2(new_n657), .A3(new_n560), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n318), .A2(new_n746), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n691), .A2(new_n751), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n741), .A2(new_n521), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n786), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n842), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n740), .A2(new_n734), .A3(new_n683), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n748), .A2(new_n850), .A3(new_n690), .A4(new_n785), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n740), .A2(new_n595), .A3(new_n664), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n775), .A3(new_n318), .A4(new_n746), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n755), .A2(new_n851), .A3(new_n853), .A4(KEYINPUT108), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n728), .A2(new_n318), .A3(new_n657), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n616), .A2(new_n736), .ZN(new_n857));
  INV_X1    g671(.A(new_n604), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n634), .A2(G472), .B1(new_n731), .B2(new_n732), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n714), .A2(new_n381), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n856), .A2(new_n613), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n614), .ZN(new_n862));
  INV_X1    g676(.A(new_n626), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n863), .A2(new_n723), .B1(new_n649), .B2(new_n659), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n469), .A2(new_n858), .A3(new_n470), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n637), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n616), .A2(new_n624), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n642), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n866), .A2(new_n868), .B1(new_n643), .B2(new_n723), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n862), .A2(new_n753), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n841), .B1(new_n855), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n724), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n649), .A2(new_n825), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n729), .A3(new_n738), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n522), .A2(new_n613), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n876), .A2(new_n658), .B1(new_n626), .B2(new_n715), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n873), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n849), .A2(new_n854), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(KEYINPUT109), .A3(new_n753), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n710), .ZN(new_n882));
  INV_X1    g696(.A(new_n743), .ZN(new_n883));
  INV_X1    g697(.A(new_n857), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n683), .A2(new_n664), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT110), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n740), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n885), .B2(new_n740), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n884), .B(new_n706), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n693), .A2(new_n882), .A3(new_n883), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT52), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n743), .B1(new_n680), .B2(new_n692), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n882), .A4(new_n889), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n892), .A2(new_n893), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT53), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n881), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n891), .A2(new_n894), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n871), .B2(new_n880), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(KEYINPUT53), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n840), .B1(new_n902), .B2(KEYINPUT54), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n897), .B(new_n900), .C1(new_n871), .C2(new_n880), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n881), .B2(new_n895), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n840), .B(KEYINPUT54), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n855), .A2(new_n870), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n895), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n910), .B(new_n911), .C1(new_n901), .C2(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n839), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n796), .B1(new_n914), .B2(new_n915), .ZN(G75));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(KEYINPUT56), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n910), .B1(new_n901), .B2(KEYINPUT53), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G902), .ZN(new_n920));
  INV_X1    g734(.A(G210), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n426), .B1(new_n430), .B2(new_n437), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n388), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT55), .Z(new_n925));
  OR2_X1    g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n925), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n266), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT117), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n926), .A2(new_n927), .A3(new_n932), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(G51));
  XNOR2_X1  g748(.A(new_n919), .B(new_n911), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n519), .B(KEYINPUT57), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n511), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n920), .A2(new_n761), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n928), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT118), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n919), .A2(G902), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n554), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n928), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT119), .Z(G60));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n913), .B2(new_n903), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n951));
  INV_X1    g765(.A(new_n621), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n950), .B2(new_n952), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n621), .A2(new_n949), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n929), .B1(new_n935), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  AND2_X1   g773(.A1(new_n919), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n654), .ZN(new_n961));
  INV_X1    g775(.A(new_n720), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n961), .B(new_n929), .C1(new_n962), .C2(new_n960), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT121), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT121), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n963), .B2(new_n965), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n603), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n596), .B1(new_n970), .B2(G224), .ZN(new_n971));
  INV_X1    g785(.A(new_n878), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n266), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n923), .B1(G898), .B2(new_n266), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  OAI22_X1  g790(.A1(new_n292), .A2(new_n293), .B1(KEYINPUT30), .B2(new_n284), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT123), .Z(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n550), .ZN(new_n979));
  INV_X1    g793(.A(new_n266), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(G900), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n768), .A2(new_n699), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n884), .A2(new_n825), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n755), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n752), .B2(new_n749), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n892), .A2(new_n882), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n779), .A2(new_n985), .A3(new_n788), .A4(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n981), .B1(new_n987), .B2(new_n980), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n707), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n868), .B(KEYINPUT125), .Z(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(new_n699), .A3(new_n747), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n788), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n993), .A2(new_n779), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n266), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n989), .B1(new_n999), .B2(new_n979), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n988), .B2(KEYINPUT126), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1000), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n998), .B2(new_n972), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n294), .A2(new_n256), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT127), .Z(new_n1008));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n283), .A3(new_n1008), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n902), .B(new_n1005), .C1(new_n703), .C2(new_n295), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n987), .B2(new_n972), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1008), .A2(new_n283), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n928), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1009), .A2(new_n1010), .A3(new_n1013), .ZN(G57));
endmodule


