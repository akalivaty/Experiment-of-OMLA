//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  OR2_X1    g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT24), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(KEYINPUT24), .B2(new_n206), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT23), .Z(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT25), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n203), .A2(KEYINPUT24), .A3(new_n204), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT25), .B1(new_n205), .B2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n210), .A2(new_n212), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n209), .B(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n212), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n204), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT28), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n214), .B(new_n218), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n226), .A2(G226gat), .A3(G233gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n226), .A2(new_n228), .B1(G226gat), .B2(G233gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231));
  INV_X1    g030(.A(G211gat), .ZN(new_n232));
  INV_X1    g031(.A(G218gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(KEYINPUT22), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G8gat), .B(G36gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G64gat), .B(G92gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n227), .B2(new_n229), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n244), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n242), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n239), .A2(KEYINPUT30), .A3(new_n243), .A4(new_n244), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n250), .A2(new_n251), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n247), .B(new_n249), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G15gat), .B(G43gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(G71gat), .B(G99gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  INV_X1    g057(.A(G227gat), .ZN(new_n259));
  INV_X1    g058(.A(G233gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT66), .B(G134gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  MUX2_X1   g063(.A(G134gat), .B(new_n264), .S(G127gat), .Z(new_n265));
  XOR2_X1   g064(.A(G113gat), .B(G120gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT67), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT68), .B(G120gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  MUX2_X1   g069(.A(G120gat), .B(new_n270), .S(G113gat), .Z(new_n271));
  XOR2_X1   g070(.A(G127gat), .B(G134gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT69), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n226), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n226), .A2(new_n276), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n262), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n258), .B1(new_n279), .B2(KEYINPUT33), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n262), .A3(new_n278), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT34), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n278), .ZN(new_n287));
  AOI221_X4 g086(.A(new_n281), .B1(KEYINPUT33), .B2(new_n258), .C1(new_n287), .C2(new_n261), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n280), .A2(new_n282), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n285), .B1(new_n291), .B2(new_n288), .ZN(new_n292));
  XOR2_X1   g091(.A(G141gat), .B(G148gat), .Z(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT2), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G155gat), .B(G162gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n228), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n237), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(G228gat), .A2(G233gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(KEYINPUT78), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(KEYINPUT78), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n308), .A2(KEYINPUT78), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n303), .A2(new_n310), .A3(new_n311), .A4(new_n306), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT79), .B(G22gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n314), .A3(new_n312), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G50gat), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT77), .B(KEYINPUT31), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n316), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(G22gat), .ZN(new_n324));
  OAI22_X1  g123(.A1(new_n316), .A2(new_n322), .B1(new_n313), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n290), .A2(new_n292), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n276), .B(new_n305), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n276), .B2(new_n305), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n305), .A2(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n276), .A3(new_n301), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n268), .A2(new_n275), .A3(KEYINPUT4), .A4(new_n299), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n329), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT74), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n337), .A2(KEYINPUT74), .A3(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G57gat), .B(G85gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT73), .B(KEYINPUT0), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT75), .B(KEYINPUT6), .Z(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n351), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n343), .B2(new_n348), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n352), .A2(KEYINPUT76), .B1(new_n355), .B2(new_n349), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n355), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n255), .B(new_n327), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n358), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT84), .B1(new_n358), .B2(KEYINPUT35), .ZN(new_n360));
  INV_X1    g159(.A(new_n326), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n290), .A2(new_n292), .A3(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n283), .A2(new_n286), .A3(KEYINPUT70), .A4(new_n289), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT35), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n348), .B(KEYINPUT81), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n343), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(new_n353), .C1(new_n348), .C2(new_n343), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n365), .A2(new_n366), .A3(new_n255), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n359), .A2(new_n360), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n330), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(KEYINPUT39), .C1(new_n330), .C2(new_n328), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(new_n367), .C1(KEYINPUT39), .C2(new_n376), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT40), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n343), .B2(new_n368), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n254), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT83), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n248), .A2(KEYINPUT37), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n248), .A2(KEYINPUT37), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n242), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT38), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n245), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(new_n389), .A3(new_n242), .A4(new_n387), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n352), .A3(new_n370), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n382), .A2(new_n254), .A3(new_n394), .A4(new_n383), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n385), .A2(new_n326), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n363), .A2(new_n364), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n397), .A2(KEYINPUT36), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT36), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n356), .A2(new_n357), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n361), .B1(new_n401), .B2(new_n254), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n202), .B1(new_n374), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n360), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n358), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n372), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(KEYINPUT85), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G43gat), .B(G50gat), .Z(new_n411));
  INV_X1    g210(.A(KEYINPUT15), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(G29gat), .A2(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT14), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT88), .B(G29gat), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n417), .A2(new_n418), .B1(G36gat), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(KEYINPUT87), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(G36gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n411), .A2(new_n412), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n414), .A2(new_n417), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(G85gat), .A3(G92gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT7), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G99gat), .A2(G106gat), .ZN(new_n432));
  INV_X1    g231(.A(G85gat), .ZN(new_n433));
  INV_X1    g232(.A(G92gat), .ZN(new_n434));
  AOI22_X1  g233(.A1(KEYINPUT8), .A2(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n428), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G99gat), .B(G106gat), .Z(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT41), .ZN(new_n440));
  NAND2_X1  g239(.A1(G232gat), .A2(G233gat), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n427), .A2(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(KEYINPUT96), .Z(new_n443));
  NAND2_X1  g242(.A1(new_n420), .A2(new_n421), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n413), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n425), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT17), .B1(new_n422), .B2(new_n426), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n439), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n441), .A2(new_n440), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT94), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n451), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G134gat), .B(G162gat), .Z(new_n455));
  XNOR2_X1  g254(.A(G190gat), .B(G218gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n457), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT16), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(G1gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(G1gat), .B2(new_n462), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n465), .A2(G8gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(G8gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469));
  NAND2_X1  g268(.A1(G71gat), .A2(G78gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G57gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(G64gat), .ZN(new_n474));
  INV_X1    g273(.A(G64gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(G57gat), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n469), .B(new_n472), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n470), .ZN(new_n478));
  NOR2_X1   g277(.A1(G71gat), .A2(G78gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n475), .A2(G57gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n473), .A2(G64gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n471), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT91), .B(new_n472), .C1(new_n474), .C2(new_n476), .ZN(new_n485));
  INV_X1    g284(.A(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT92), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n468), .B1(new_n492), .B2(KEYINPUT21), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(new_n232), .ZN(new_n494));
  XOR2_X1   g293(.A(G127gat), .B(G155gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n492), .A2(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g296(.A1(G231gat), .A2(G233gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n496), .B(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT93), .B(G183gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n500), .B(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n461), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n438), .A2(KEYINPUT98), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n437), .B(new_n509), .Z(new_n510));
  INV_X1    g309(.A(new_n488), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n484), .A2(KEYINPUT92), .A3(new_n487), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT92), .B1(new_n484), .B2(new_n487), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT97), .B1(new_n516), .B2(new_n439), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n490), .A2(KEYINPUT97), .A3(new_n439), .A4(new_n491), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n508), .B(new_n513), .C1(new_n517), .C2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n439), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n492), .A2(KEYINPUT10), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n507), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n490), .A2(new_n491), .A3(new_n439), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n512), .B1(new_n527), .B2(new_n518), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(new_n506), .ZN(new_n529));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G176gat), .B(G204gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n524), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n535));
  INV_X1    g334(.A(new_n522), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n528), .B2(new_n508), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n537), .B2(new_n507), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n522), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT99), .A3(new_n506), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n540), .A3(new_n529), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n534), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n410), .A2(new_n505), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n468), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT90), .B1(new_n427), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n445), .A2(new_n425), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n468), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n547), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT89), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT13), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n449), .A2(new_n544), .ZN(new_n556));
  INV_X1    g355(.A(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n547), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n557), .A4(new_n547), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT86), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  INV_X1    g364(.A(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT11), .B(G169gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT12), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n562), .A2(new_n563), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n543), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n401), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g378(.A1(new_n543), .A2(new_n575), .A3(new_n254), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G8gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT42), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n580), .A2(KEYINPUT42), .A3(new_n583), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT101), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n580), .A2(new_n588), .A3(G8gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n580), .B2(G8gat), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n586), .A2(new_n587), .B1(new_n590), .B2(new_n591), .ZN(G1325gat));
  INV_X1    g391(.A(G15gat), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n576), .A2(new_n593), .A3(new_n400), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n543), .A2(new_n575), .A3(new_n397), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(G1326gat));
  NOR2_X1   g395(.A1(new_n576), .A2(new_n326), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT43), .B(G22gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(G1327gat));
  INV_X1    g398(.A(new_n504), .ZN(new_n600));
  INV_X1    g399(.A(new_n542), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n600), .A2(new_n574), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n410), .A2(new_n461), .A3(new_n602), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n603), .A2(new_n577), .A3(new_n419), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT45), .Z(new_n605));
  INV_X1    g404(.A(new_n419), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n404), .A2(new_n461), .A3(new_n409), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT44), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n374), .B2(new_n403), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n407), .A2(KEYINPUT102), .A3(new_n408), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n460), .A2(KEYINPUT44), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n615), .A2(new_n602), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n616), .A2(new_n401), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n605), .B1(new_n606), .B2(new_n617), .ZN(G1328gat));
  NOR3_X1   g417(.A1(new_n603), .A2(G36gat), .A3(new_n255), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT46), .ZN(new_n620));
  INV_X1    g419(.A(G36gat), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n616), .A2(new_n254), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(G1329gat));
  INV_X1    g422(.A(new_n400), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n616), .A2(G43gat), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G43gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n397), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n603), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT47), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT47), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n625), .A2(new_n631), .A3(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(G1330gat));
  NAND3_X1  g432(.A1(new_n615), .A2(new_n361), .A3(new_n602), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n615), .A2(new_n636), .A3(new_n361), .A4(new_n602), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(G50gat), .A3(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n603), .A2(G50gat), .A3(new_n326), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(KEYINPUT48), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT48), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n634), .A2(G50gat), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(G1331gat));
  AND2_X1   g444(.A1(new_n612), .A2(new_n505), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n575), .A2(new_n542), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n577), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(new_n473), .ZN(G1332gat));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n255), .ZN(new_n651));
  NOR2_X1   g450(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n652));
  AND2_X1   g451(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n651), .B2(new_n652), .ZN(G1333gat));
  NAND4_X1  g454(.A1(new_n646), .A2(G71gat), .A3(new_n624), .A4(new_n647), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n648), .A2(new_n627), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(G71gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1334gat));
  NOR2_X1   g459(.A1(new_n648), .A2(new_n326), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(G78gat), .Z(G1335gat));
  NAND3_X1  g461(.A1(new_n615), .A2(new_n504), .A3(new_n647), .ZN(new_n663));
  OAI21_X1  g462(.A(G85gat), .B1(new_n663), .B2(new_n577), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n460), .A2(new_n575), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n504), .B(new_n665), .C1(new_n374), .C2(new_n403), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT51), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT105), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n433), .A3(new_n601), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n664), .B1(new_n670), .B2(new_n577), .ZN(G1336gat));
  NAND4_X1  g470(.A1(new_n668), .A2(new_n434), .A3(new_n601), .A4(new_n254), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT106), .B(KEYINPUT52), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n607), .A2(KEYINPUT44), .B1(new_n612), .B2(new_n613), .ZN(new_n674));
  INV_X1    g473(.A(new_n647), .ZN(new_n675));
  NOR4_X1   g474(.A1(new_n674), .A2(new_n600), .A3(new_n255), .A4(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n672), .B(new_n673), .C1(new_n676), .C2(new_n434), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT107), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n674), .A2(new_n600), .A3(new_n675), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n434), .B1(new_n679), .B2(new_n254), .ZN(new_n680));
  INV_X1    g479(.A(new_n672), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT52), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G92gat), .B1(new_n663), .B2(new_n255), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n672), .A4(new_n673), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n678), .A2(new_n682), .A3(new_n685), .ZN(G1337gat));
  XOR2_X1   g485(.A(KEYINPUT108), .B(G99gat), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n601), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n663), .A2(new_n400), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n688), .A2(new_n627), .B1(new_n689), .B2(new_n687), .ZN(G1338gat));
  NAND2_X1  g489(.A1(new_n668), .A2(new_n601), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(G106gat), .A3(new_n326), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n663), .A2(new_n326), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT109), .B(G106gat), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n694), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n679), .B2(new_n361), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(new_n692), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(G1339gat));
  INV_X1    g500(.A(new_n534), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n538), .B2(new_n540), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n520), .A2(new_n507), .A3(new_n522), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT54), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n532), .B1(new_n707), .B2(new_n523), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT112), .B1(new_n709), .B2(KEYINPUT55), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT99), .B1(new_n539), .B2(new_n506), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n535), .B(new_n507), .C1(new_n520), .C2(new_n522), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n703), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT54), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n537), .B2(new_n507), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n533), .B1(new_n715), .B2(new_n524), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n713), .A2(new_n716), .A3(KEYINPUT112), .A4(KEYINPUT55), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n702), .B1(new_n710), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT113), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n713), .A2(new_n716), .A3(KEYINPUT55), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n717), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n702), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n571), .B(new_n573), .C1(KEYINPUT55), .C2(new_n709), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n720), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n562), .A2(new_n570), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n550), .A2(new_n554), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n557), .B1(new_n556), .B2(new_n547), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n730), .B1(new_n569), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n601), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n729), .A2(KEYINPUT114), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT114), .B1(new_n729), .B2(new_n735), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n736), .A2(new_n737), .A3(new_n461), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739));
  INV_X1    g538(.A(new_n709), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n460), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n741), .A2(new_n734), .A3(new_n720), .A4(new_n726), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n504), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NOR4_X1   g543(.A1(new_n461), .A2(new_n504), .A3(new_n575), .A4(new_n601), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n401), .A3(new_n327), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n254), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n574), .A2(G113gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT116), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n747), .A2(new_n401), .A3(new_n255), .A4(new_n365), .ZN(new_n755));
  OAI21_X1  g554(.A(G113gat), .B1(new_n755), .B2(new_n574), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1340gat));
  NAND3_X1  g556(.A1(new_n751), .A2(new_n270), .A3(new_n601), .ZN(new_n758));
  OAI21_X1  g557(.A(G120gat), .B1(new_n755), .B2(new_n542), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1341gat));
  NOR3_X1   g559(.A1(new_n748), .A2(new_n504), .A3(new_n254), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n600), .A2(G127gat), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n761), .A2(G127gat), .B1(new_n755), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT117), .Z(G1342gat));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n264), .A3(new_n461), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n765), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT56), .ZN(new_n767));
  OAI21_X1  g566(.A(G134gat), .B1(new_n755), .B2(new_n460), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT118), .B1(new_n765), .B2(KEYINPUT56), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(G1343gat));
  AOI21_X1  g569(.A(new_n326), .B1(new_n744), .B2(new_n746), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT120), .B1(new_n771), .B2(KEYINPUT57), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n735), .B1(new_n719), .B2(new_n727), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n735), .B(KEYINPUT121), .C1(new_n719), .C2(new_n727), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n460), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n600), .B1(new_n777), .B2(new_n742), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n361), .B1(new_n778), .B2(new_n745), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n725), .B1(new_n724), .B2(new_n702), .ZN(new_n784));
  AOI211_X1 g583(.A(KEYINPUT113), .B(new_n534), .C1(new_n723), .C2(new_n717), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n784), .A2(new_n785), .A3(new_n727), .ZN(new_n786));
  INV_X1    g585(.A(new_n735), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n729), .A2(KEYINPUT114), .A3(new_n735), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n460), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n600), .B1(new_n790), .B2(new_n742), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n745), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n782), .B(new_n780), .C1(new_n792), .C2(new_n326), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n772), .A2(new_n781), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n624), .A2(new_n577), .A3(new_n254), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT119), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n794), .A2(G141gat), .A3(new_n575), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(G141gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n771), .A2(new_n795), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n574), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(KEYINPUT58), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1344gat));
  NAND3_X1  g605(.A1(new_n794), .A2(new_n601), .A3(new_n797), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(G148gat), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n361), .C1(new_n791), .C2(new_n745), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n779), .A2(new_n780), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n601), .ZN(new_n813));
  OAI21_X1  g612(.A(G148gat), .B1(new_n813), .B2(new_n796), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT59), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n800), .A2(G148gat), .A3(new_n542), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT122), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1345gat));
  NAND4_X1  g618(.A1(new_n794), .A2(G155gat), .A3(new_n600), .A4(new_n797), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n294), .B1(new_n800), .B2(new_n504), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(G1346gat));
  NAND3_X1  g621(.A1(new_n794), .A2(new_n461), .A3(new_n797), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n794), .A2(KEYINPUT123), .A3(new_n461), .A4(new_n797), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(G162gat), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n771), .A2(new_n295), .A3(new_n461), .A4(new_n795), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1347gat));
  NAND4_X1  g628(.A1(new_n747), .A2(new_n577), .A3(new_n254), .A4(new_n365), .ZN(new_n830));
  OAI21_X1  g629(.A(G169gat), .B1(new_n830), .B2(new_n574), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n747), .A2(new_n577), .A3(new_n254), .A4(new_n327), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(G169gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n833), .B2(new_n574), .ZN(G1348gat));
  INV_X1    g633(.A(new_n832), .ZN(new_n835));
  AOI21_X1  g634(.A(G176gat), .B1(new_n835), .B2(new_n601), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n830), .A2(new_n542), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(G176gat), .B2(new_n837), .ZN(G1349gat));
  OAI21_X1  g637(.A(G183gat), .B1(new_n830), .B2(new_n504), .ZN(new_n839));
  INV_X1    g638(.A(new_n222), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT124), .B1(new_n841), .B2(new_n600), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n832), .A2(new_n843), .A3(new_n504), .A4(new_n840), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT60), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n839), .B(new_n847), .C1(new_n842), .C2(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1350gat));
  OAI21_X1  g648(.A(G190gat), .B1(new_n830), .B2(new_n460), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n223), .A3(new_n461), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1351gat));
  NAND3_X1  g654(.A1(new_n400), .A2(new_n577), .A3(new_n254), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n810), .B2(new_n811), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n566), .B1(new_n857), .B2(new_n575), .ZN(new_n858));
  INV_X1    g657(.A(new_n856), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n771), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(G197gat), .A3(new_n574), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n858), .A2(new_n861), .ZN(G1352gat));
  NOR3_X1   g661(.A1(new_n860), .A2(G204gat), .A3(new_n542), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G204gat), .B1(new_n813), .B2(new_n856), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n864), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1353gat));
  NAND4_X1  g667(.A1(new_n771), .A2(new_n232), .A3(new_n600), .A4(new_n859), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(new_n232), .C1(new_n857), .C2(new_n600), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n812), .A2(new_n600), .A3(new_n859), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT63), .B1(new_n872), .B2(G211gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT126), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n869), .C1(new_n871), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1354gat));
  NAND2_X1  g677(.A1(new_n812), .A2(new_n859), .ZN(new_n879));
  OAI21_X1  g678(.A(G218gat), .B1(new_n879), .B2(new_n460), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n461), .A2(new_n233), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n860), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


