//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n207), .A2(G13), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  AND2_X1   g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n218), .B(new_n222), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n232), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n246), .A2(G222), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n246), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n248), .B1(new_n249), .B2(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n223), .B2(new_n253), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n255), .A2(new_n261), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(G226), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G179), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  INV_X1    g0075(.A(new_n273), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n271), .ZN(new_n277));
  OR3_X1    g0077(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT67), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n259), .A2(G20), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  OAI21_X1  g0081(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n282), .B1(new_n283), .B2(new_n285), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(new_n277), .B1(new_n290), .B2(new_n276), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n269), .B(new_n292), .C1(G169), .C2(new_n267), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n292), .B(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n266), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(G200), .B2(new_n266), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n294), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n276), .A2(new_n209), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n284), .A2(G50), .B1(G20), .B2(new_n209), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n249), .B2(new_n288), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT11), .A3(new_n277), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n279), .A2(G68), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n305), .B(new_n308), .C1(new_n274), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT11), .B1(new_n307), .B2(new_n277), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n263), .B1(G238), .B2(new_n264), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n246), .A2(G226), .A3(new_n247), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n323), .A2(new_n234), .A3(new_n247), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n255), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n315), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n315), .B2(new_n325), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n314), .B(G169), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n329), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n327), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n268), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n314), .B1(new_n332), .B2(G169), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n313), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(G200), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(new_n312), .C1(new_n296), .C2(new_n332), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G20), .A2(G77), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n338), .B1(new_n286), .B2(new_n285), .C1(new_n288), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n277), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n279), .A2(G77), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(G77), .B2(new_n273), .C1(new_n274), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G107), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n250), .A2(new_n210), .B1(new_n344), .B2(new_n246), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n323), .A2(new_n234), .A3(G1698), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n255), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n263), .B1(G244), .B2(new_n264), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n343), .B1(G190), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n350), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G169), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n343), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n349), .A2(G179), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n303), .A2(new_n335), .A3(new_n337), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n254), .A2(G232), .A3(new_n260), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n254), .A2(new_n260), .A3(KEYINPUT69), .A4(G232), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n262), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT70), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n364), .A2(KEYINPUT70), .A3(new_n262), .A4(new_n365), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n320), .A2(new_n322), .A3(G226), .A4(G1698), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n320), .A2(new_n322), .A3(G223), .A4(new_n247), .ZN(new_n371));
  AND3_X1   g0171(.A1(KEYINPUT68), .A2(G33), .A3(G87), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT68), .B1(G33), .B2(G87), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(G190), .B1(new_n375), .B2(new_n255), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n368), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n375), .A2(new_n255), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n352), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n323), .B2(new_n287), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n382), .B(G20), .C1(new_n320), .C2(new_n322), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n284), .A2(G159), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n209), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n201), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n382), .B1(new_n246), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n323), .A2(KEYINPUT7), .A3(new_n287), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n209), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n385), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n389), .A2(new_n395), .A3(new_n277), .ZN(new_n396));
  INV_X1    g0196(.A(new_n286), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n273), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n280), .B2(new_n397), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n380), .A2(KEYINPUT72), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n380), .A2(KEYINPUT71), .A3(new_n396), .A4(new_n399), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT17), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n403), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n368), .A2(new_n369), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n378), .A2(G179), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n378), .A2(new_n366), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n409), .A2(new_n410), .B1(new_n411), .B2(new_n355), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n396), .A2(new_n399), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT18), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n361), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G283), .ZN(new_n421));
  INV_X1    g0221(.A(G97), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n287), .C1(G33), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G116), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G20), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n277), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n270), .A2(new_n271), .B1(G20), .B2(new_n424), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(KEYINPUT20), .A3(new_n423), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n273), .A2(G116), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n259), .A2(G33), .ZN(new_n433));
  AND4_X1   g0233(.A1(new_n271), .A2(new_n273), .A3(new_n270), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n434), .B2(G116), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n355), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n321), .A2(G33), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n438));
  OAI21_X1  g0238(.A(G303), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n320), .A2(new_n322), .A3(G264), .A4(G1698), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n320), .A2(new_n322), .A3(G257), .A4(new_n247), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n255), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT5), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(G41), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G270), .A3(new_n254), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n258), .A2(new_n446), .A3(new_n448), .A4(new_n450), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n451), .A2(KEYINPUT79), .A3(G270), .A4(new_n254), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n443), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n436), .A2(new_n457), .A3(KEYINPUT21), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n268), .B1(new_n431), .B2(new_n435), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n454), .A2(new_n456), .ZN(new_n460));
  INV_X1    g0260(.A(new_n455), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n442), .B2(new_n255), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n457), .A2(G200), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n429), .A2(KEYINPUT20), .A3(new_n423), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n429), .B2(new_n423), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n432), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n272), .A2(new_n273), .A3(new_n433), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n424), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n465), .B(new_n472), .C1(new_n296), .C2(new_n457), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n436), .A2(new_n457), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(KEYINPUT80), .B(KEYINPUT21), .C1(new_n436), .C2(new_n457), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n464), .B(new_n473), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n480));
  AND4_X1   g0280(.A1(new_n443), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n481));
  OAI21_X1  g0281(.A(G169), .B1(new_n468), .B2(new_n471), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n475), .A2(new_n474), .A3(new_n476), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n464), .A4(new_n473), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G107), .B1(new_n381), .B2(new_n383), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  AND2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n204), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n344), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n272), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n273), .A2(G97), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n434), .B2(G97), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n497), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n284), .A2(G77), .ZN(new_n503));
  INV_X1    g0303(.A(new_n494), .ZN(new_n504));
  XNOR2_X1  g0304(.A(G97), .B(G107), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n491), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n503), .B1(new_n506), .B2(new_n287), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n344), .B1(new_n391), .B2(new_n392), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n277), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n509), .B2(new_n499), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n320), .A2(new_n322), .A3(G244), .A4(new_n247), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G250), .A2(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT4), .A2(G244), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G1698), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n246), .A2(new_n517), .B1(G33), .B2(G283), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n254), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n451), .A2(G257), .A3(new_n254), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n455), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT75), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT75), .B1(new_n519), .B2(new_n521), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(KEYINPUT76), .A3(G200), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT76), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(G200), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n519), .A2(new_n521), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G190), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n511), .A2(new_n525), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n514), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n255), .ZN(new_n533));
  INV_X1    g0333(.A(new_n521), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G169), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n529), .A2(G179), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n497), .B2(new_n500), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n258), .A2(new_n448), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n254), .B(G250), .C1(G1), .C2(new_n447), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n320), .A2(new_n322), .A3(G244), .A4(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT77), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT77), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n246), .A2(new_n546), .A3(G244), .A4(G1698), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n246), .A2(G238), .A3(new_n247), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n543), .B1(new_n550), .B2(new_n255), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(G169), .ZN(new_n552));
  AOI211_X1 g0352(.A(G179), .B(new_n543), .C1(new_n550), .C2(new_n255), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n287), .B1(new_n317), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G87), .B2(new_n205), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n320), .A2(new_n322), .A3(new_n287), .A4(G68), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n555), .B1(new_n288), .B2(new_n422), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n277), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n339), .A2(new_n276), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n470), .A2(new_n339), .ZN(new_n563));
  AND4_X1   g0363(.A1(KEYINPUT78), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n560), .A2(new_n277), .B1(new_n276), .B2(new_n339), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT78), .B1(new_n565), .B2(new_n563), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n551), .A2(new_n352), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n434), .A2(G87), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n561), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(G190), .B2(new_n551), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n554), .A2(new_n567), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n451), .A2(G264), .A3(new_n254), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT83), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n451), .A2(new_n575), .A3(G264), .A4(new_n254), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n320), .A2(new_n322), .A3(G257), .A4(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n320), .A2(new_n322), .A3(G250), .A4(new_n247), .ZN(new_n579));
  INV_X1    g0379(.A(G294), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n579), .C1(new_n319), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n255), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n455), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n352), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n461), .B1(new_n574), .B2(new_n576), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(KEYINPUT82), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT82), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n587), .A3(new_n255), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n584), .B1(G190), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n320), .A2(new_n322), .A3(new_n287), .A4(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT22), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n246), .A2(new_n593), .A3(new_n287), .A4(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n548), .A2(G20), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT23), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n287), .B2(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n344), .A2(KEYINPUT23), .A3(G20), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n272), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT25), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n273), .B2(G107), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n273), .A2(new_n606), .A3(G107), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n344), .A2(new_n470), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n590), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n581), .A2(new_n587), .A3(new_n255), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n587), .B1(new_n581), .B2(new_n255), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n355), .B1(new_n615), .B2(new_n585), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n585), .A2(G179), .A3(new_n582), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n616), .A2(new_n618), .B1(new_n605), .B2(new_n610), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n572), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n540), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n420), .A2(new_n489), .A3(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n551), .A2(new_n268), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n565), .A2(new_n563), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n550), .A2(new_n255), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT84), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n550), .A2(KEYINPUT84), .A3(new_n255), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n543), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n623), .B(new_n624), .C1(new_n629), .C2(G169), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n486), .A2(new_n464), .A3(new_n619), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n539), .A3(new_n531), .A4(new_n612), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n623), .A2(new_n624), .ZN(new_n633));
  INV_X1    g0433(.A(new_n543), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n550), .A2(KEYINPUT84), .A3(new_n255), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT84), .B1(new_n550), .B2(new_n255), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n355), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n625), .A2(G190), .A3(new_n634), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n561), .A2(new_n562), .A3(new_n569), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(G200), .B2(new_n637), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT85), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n638), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n571), .B1(new_n629), .B2(new_n352), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT85), .B1(new_n630), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n630), .B1(new_n632), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n539), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n572), .A3(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n643), .B1(new_n638), .B2(new_n642), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n630), .A2(KEYINPUT85), .A3(new_n645), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n538), .B1(new_n501), .B2(new_n510), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n651), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n420), .B1(new_n648), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n418), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n337), .A2(new_n359), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n335), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n407), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n300), .A2(new_n302), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n294), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n259), .A2(new_n287), .A3(G13), .ZN(new_n668));
  OAI21_X1  g0468(.A(G213), .B1(new_n668), .B2(KEYINPUT27), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(KEYINPUT27), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n472), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n480), .B2(new_n488), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n673), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n612), .A2(new_n619), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n611), .B2(new_n672), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n619), .B2(new_n672), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n672), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n486), .B2(new_n464), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n619), .B2(new_n684), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n683), .A2(new_n687), .ZN(G399));
  NAND2_X1  g0488(.A1(new_n220), .A2(new_n449), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT87), .B1(new_n690), .B2(new_n227), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(G1), .A3(new_n692), .ZN(new_n693));
  MUX2_X1   g0493(.A(KEYINPUT87), .B(new_n691), .S(new_n693), .Z(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT26), .B1(new_n649), .B2(new_n572), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n655), .B1(new_n652), .B2(new_n653), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(KEYINPUT26), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT29), .B(new_n672), .C1(new_n648), .C2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n531), .A2(new_n539), .A3(new_n612), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n589), .A2(G169), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n602), .A2(new_n604), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n277), .ZN(new_n704));
  INV_X1    g0504(.A(new_n610), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n617), .A2(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n675), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n638), .B1(new_n708), .B2(new_n654), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n650), .B1(new_n698), .B2(KEYINPUT26), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n684), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n700), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT90), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n577), .A2(new_n582), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n457), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n535), .A2(new_n268), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT30), .A4(new_n551), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n460), .A2(new_n462), .A3(new_n577), .A4(new_n582), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n551), .A2(new_n529), .A3(G179), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n481), .A2(G179), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n583), .A2(KEYINPUT89), .A3(new_n535), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT89), .B1(new_n583), .B2(new_n535), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n637), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n714), .B(new_n672), .C1(new_n723), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n722), .A3(new_n718), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n729), .B2(new_n684), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n621), .A2(new_n489), .A3(new_n672), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n712), .A2(new_n713), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n713), .B1(new_n712), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n696), .B1(new_n738), .B2(G1), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT91), .ZN(G364));
  INV_X1    g0540(.A(new_n678), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n676), .A2(new_n677), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n287), .A2(G13), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n259), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n690), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n741), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n676), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n220), .A2(new_n323), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT92), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n244), .A2(G45), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(G45), .C2(new_n226), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n220), .A2(new_n246), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n756), .B1(G116), .B2(new_n220), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n271), .B1(G20), .B2(new_n355), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n751), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n747), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n760), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n287), .A2(new_n296), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n352), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n323), .B1(new_n767), .B2(G87), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n296), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n287), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n287), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n765), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n768), .B1(new_n422), .B2(new_n770), .C1(new_n344), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n771), .A2(new_n268), .A3(new_n352), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT95), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n781));
  XNOR2_X1  g0581(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n287), .A2(new_n268), .A3(new_n352), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n783), .A2(KEYINPUT97), .A3(new_n296), .ZN(new_n784));
  AOI21_X1  g0584(.A(KEYINPUT97), .B1(new_n783), .B2(new_n296), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n773), .B(new_n782), .C1(G68), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n783), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n296), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n764), .A2(G179), .A3(new_n352), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n290), .B1(new_n386), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n771), .A2(G179), .A3(new_n352), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n795), .A2(KEYINPUT93), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(KEYINPUT93), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n793), .B1(new_n799), .B2(G77), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT94), .Z(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n770), .A2(new_n580), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G326), .B2(new_n790), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  NOR2_X1   g0606(.A1(new_n786), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n792), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G322), .B1(new_n767), .B2(G303), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n323), .C1(new_n810), .C2(new_n772), .ZN(new_n811));
  INV_X1    g0611(.A(new_n778), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n807), .B(new_n811), .C1(G329), .C2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n788), .A2(new_n801), .B1(new_n805), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n752), .B(new_n762), .C1(new_n763), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n748), .A2(new_n815), .ZN(G396));
  AOI22_X1  g0616(.A1(new_n799), .A2(G116), .B1(G311), .B2(new_n812), .ZN(new_n817));
  INV_X1    g0617(.A(G303), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n791), .A2(new_n818), .B1(new_n770), .B2(new_n422), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n323), .B1(new_n792), .B2(new_n580), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n766), .A2(new_n344), .B1(new_n772), .B2(new_n211), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n817), .B(new_n822), .C1(new_n810), .C2(new_n786), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n790), .A2(G137), .B1(G143), .B2(new_n808), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n283), .B2(new_n786), .C1(new_n798), .C2(new_n779), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  OAI21_X1  g0626(.A(new_n246), .B1(new_n772), .B2(new_n209), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G50), .B2(new_n767), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n386), .B2(new_n770), .C1(new_n829), .C2(new_n778), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT100), .Z(new_n831));
  OAI21_X1  g0631(.A(new_n823), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n760), .A2(new_n749), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n832), .A2(new_n760), .B1(new_n249), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT101), .B1(new_n357), .B2(new_n358), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n684), .A2(new_n343), .ZN(new_n838));
  INV_X1    g0638(.A(new_n358), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT101), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n343), .A4(new_n356), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n353), .A2(new_n837), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n359), .A2(new_n684), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n836), .B1(new_n845), .B2(new_n750), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n746), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n844), .B(KEYINPUT102), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(new_n711), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n837), .A2(new_n841), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n353), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n672), .B(new_n852), .C1(new_n659), .C2(new_n648), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n849), .A2(new_n734), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n747), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n734), .B1(new_n849), .B2(new_n853), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n847), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT103), .Z(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  OR2_X1    g0659(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(G116), .A4(new_n225), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT36), .Z(new_n863));
  OR3_X1    g0663(.A1(new_n226), .A2(new_n249), .A3(new_n387), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n290), .A2(G68), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n259), .B(G13), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT106), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n733), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT106), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n335), .A2(new_n872), .A3(new_n337), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n313), .A2(new_n684), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n335), .A2(KEYINPUT104), .A3(new_n337), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n333), .A2(new_n334), .A3(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n845), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n413), .A2(new_n670), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT105), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT105), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n413), .A2(new_n884), .A3(new_n670), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n407), .B2(new_n418), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n380), .A2(new_n396), .A3(new_n399), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n414), .A2(new_n888), .A3(new_n889), .A4(new_n882), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n396), .A2(new_n399), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n355), .B1(new_n378), .B2(new_n366), .ZN(new_n892));
  INV_X1    g0692(.A(new_n410), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n408), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n889), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n883), .B2(new_n885), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n890), .B1(new_n896), .B2(new_n888), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n887), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT40), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n881), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n882), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n407), .B2(new_n418), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n895), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n890), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n901), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(new_n869), .A3(new_n870), .A4(new_n879), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n871), .A2(new_n419), .A3(new_n361), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n913), .A2(new_n914), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n916), .A2(new_n917), .A3(new_n677), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n875), .A2(new_n878), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n850), .A2(new_n684), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n853), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n900), .A2(new_n901), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n887), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n908), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n335), .A2(new_n684), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n661), .A2(new_n670), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n924), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n420), .B(new_n700), .C1(new_n711), .C2(KEYINPUT29), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n666), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n918), .A2(new_n937), .B1(new_n259), .B2(new_n743), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n918), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n867), .B1(new_n938), .B2(new_n939), .ZN(G367));
  AND2_X1   g0740(.A1(new_n754), .A2(new_n231), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n761), .B1(new_n220), .B2(new_n339), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n746), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n770), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n790), .A2(G143), .B1(new_n944), .B2(G68), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n323), .B1(new_n767), .B2(G58), .ZN(new_n946));
  INV_X1    g0746(.A(new_n772), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n808), .A2(G150), .B1(new_n947), .B2(G77), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(G137), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n798), .A2(new_n290), .B1(new_n950), .B2(new_n778), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n949), .B(new_n951), .C1(G159), .C2(new_n787), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT110), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n323), .B1(new_n772), .B2(new_n422), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G303), .B2(new_n808), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n955), .B1(new_n956), .B2(new_n778), .C1(new_n798), .C2(new_n810), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n766), .A2(new_n424), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT46), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G311), .B2(new_n790), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G107), .A2(new_n944), .B1(new_n958), .B2(KEYINPUT46), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n580), .C2(new_n786), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n953), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n943), .B1(new_n964), .B2(new_n760), .ZN(new_n965));
  INV_X1    g0765(.A(new_n751), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n654), .B1(new_n640), .B2(new_n672), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n638), .A2(new_n570), .A3(new_n684), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n511), .A2(new_n672), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n540), .A2(new_n971), .B1(new_n655), .B2(new_n672), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT108), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(new_n686), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT42), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n539), .B1(new_n973), .B2(new_n619), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n672), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n969), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n981), .B2(new_n979), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n975), .B2(new_n977), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n682), .A2(new_n973), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n973), .A2(new_n687), .ZN(new_n992));
  NOR2_X1   g0792(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n973), .A2(new_n687), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n683), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n999), .A3(new_n682), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n686), .B1(new_n681), .B2(new_n685), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n678), .B(new_n1004), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n738), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n689), .B(KEYINPUT41), .Z(new_n1007));
  AOI21_X1  g0807(.A(new_n745), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n970), .B1(new_n991), .B2(new_n1008), .ZN(G387));
  NOR2_X1   g0809(.A1(new_n737), .A2(new_n1005), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n737), .A2(new_n1005), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n690), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1005), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n681), .A2(new_n966), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n758), .A2(new_n692), .B1(G107), .B2(new_n220), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n754), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n692), .B(new_n447), .C1(new_n209), .C2(new_n249), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT50), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n286), .B2(G50), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n397), .A2(KEYINPUT50), .A3(new_n290), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1017), .A2(KEYINPUT111), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G45), .B2(new_n237), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT111), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1016), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n761), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n746), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n246), .B1(new_n772), .B2(new_n422), .C1(new_n770), .C2(new_n339), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n767), .A2(G77), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n290), .B2(new_n792), .C1(new_n209), .C2(new_n794), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(new_n397), .C2(new_n787), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT112), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n791), .B2(new_n779), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n790), .A2(KEYINPUT112), .A3(G159), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n812), .A2(G150), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n812), .A2(G326), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n246), .B1(new_n947), .B2(G116), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n770), .A2(new_n810), .B1(new_n766), .B2(new_n580), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n790), .A2(G322), .B1(G317), .B2(new_n808), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n802), .B2(new_n786), .C1(new_n798), .C2(new_n818), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1038), .B(new_n1039), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1028), .B1(new_n1049), .B2(new_n760), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1014), .A2(new_n745), .B1(new_n1015), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1013), .A2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1003), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n1010), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1055), .A3(new_n690), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n973), .A2(new_n751), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n754), .A2(new_n241), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n761), .B1(new_n220), .B2(new_n422), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n746), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n799), .A2(new_n397), .B1(G143), .B2(new_n812), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n246), .B1(new_n772), .B2(new_n211), .C1(new_n209), .C2(new_n766), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G77), .B2(new_n944), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n290), .C2(new_n786), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n790), .A2(G150), .B1(G159), .B2(new_n808), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n580), .A2(new_n794), .B1(new_n766), .B2(new_n810), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n246), .B(new_n1067), .C1(G107), .C2(new_n947), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n787), .A2(G303), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n812), .A2(G322), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n944), .A2(G116), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n790), .A2(G317), .B1(G311), .B2(new_n808), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1064), .A2(new_n1066), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1060), .B1(new_n1075), .B2(new_n760), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1054), .A2(new_n745), .B1(new_n1057), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1056), .A2(new_n1077), .ZN(G390));
  NAND4_X1  g0878(.A1(new_n869), .A2(new_n879), .A3(G330), .A4(new_n870), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n927), .A2(new_n928), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n922), .B2(new_n930), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n672), .B(new_n852), .C1(new_n648), .C2(new_n699), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n921), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n919), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n930), .B1(new_n909), .B2(new_n901), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1079), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT113), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n684), .B(new_n851), .C1(new_n709), .C2(new_n710), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1090), .B2(new_n920), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1091), .A2(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n910), .A2(new_n929), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n919), .B1(new_n1082), .B2(new_n921), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n733), .A2(G330), .A3(new_n845), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1093), .A2(new_n1094), .B1(new_n919), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n919), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n1081), .A3(KEYINPUT113), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1088), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1080), .A2(new_n749), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n746), .B1(new_n834), .B2(new_n397), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n799), .A2(G97), .B1(G294), .B2(new_n812), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n792), .A2(new_n424), .B1(new_n772), .B2(new_n209), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n246), .B(new_n1105), .C1(G87), .C2(new_n767), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n790), .A2(G283), .B1(new_n944), .B2(G77), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n786), .A2(new_n344), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n246), .B1(new_n792), .B2(new_n829), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G50), .B2(new_n947), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n778), .C1(new_n798), .C2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n766), .A2(new_n283), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n790), .A2(G128), .B1(new_n944), .B2(G159), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n950), .C2(new_n786), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1108), .A2(new_n1109), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1120), .B2(new_n760), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1101), .A2(new_n745), .B1(new_n1102), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n869), .A2(new_n420), .A3(G330), .A4(new_n870), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n934), .A2(new_n1123), .A3(new_n666), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n677), .B(new_n844), .C1(new_n731), .C2(new_n732), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT114), .B1(new_n1125), .B2(new_n1084), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT114), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1095), .A2(new_n1127), .A3(new_n919), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1079), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n853), .A2(new_n921), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1098), .A2(new_n1083), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n869), .A2(new_n848), .A3(G330), .A4(new_n870), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n919), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1124), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n690), .B1(new_n1101), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1079), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT113), .B1(new_n1099), .B2(new_n1081), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1099), .A2(new_n1081), .A3(KEYINPUT113), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1136), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1122), .B1(new_n1137), .B2(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT118), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1147), .B(new_n1124), .C1(new_n1101), .C2(new_n1136), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1124), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT118), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n881), .A2(new_n902), .B1(new_n911), .B2(KEYINPUT40), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n292), .A2(new_n670), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n303), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n303), .A2(new_n1153), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1152), .A2(new_n677), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1161), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n913), .B2(G330), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n933), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1161), .B1(new_n1152), .B2(new_n677), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n913), .A2(G330), .A3(new_n1163), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n933), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1146), .B1(new_n1151), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1146), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n690), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(new_n745), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1161), .A2(new_n749), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n747), .B1(new_n290), .B2(new_n833), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT116), .Z(new_n1179));
  NOR2_X1   g0979(.A1(new_n246), .A2(G41), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G50), .B(new_n1180), .C1(new_n319), .C2(new_n449), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n947), .A2(G58), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n344), .B2(new_n792), .C1(new_n339), .C2(new_n794), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G283), .B2(new_n812), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1030), .B(new_n1180), .C1(new_n209), .C2(new_n770), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G116), .B2(new_n790), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(new_n422), .C2(new_n786), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT58), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1181), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(G128), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n792), .A2(new_n1190), .B1(new_n766), .B2(new_n1113), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G137), .B2(new_n795), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n790), .A2(G125), .B1(new_n944), .B2(G150), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n829), .C2(new_n786), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n812), .A2(G124), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n947), .C2(G159), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1189), .B1(new_n1188), .B2(new_n1187), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1179), .B1(new_n1200), .B2(new_n760), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1177), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1176), .A2(KEYINPUT117), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT117), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n744), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1202), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1175), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(G375));
  AOI22_X1  g1010(.A1(new_n799), .A2(G107), .B1(G303), .B2(new_n812), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n791), .A2(new_n580), .B1(new_n770), .B2(new_n339), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n323), .B1(new_n772), .B2(new_n249), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n792), .A2(new_n810), .B1(new_n766), .B2(new_n422), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1211), .B(new_n1215), .C1(new_n424), .C2(new_n786), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n786), .A2(new_n1113), .ZN(new_n1217));
  OR3_X1    g1017(.A1(new_n791), .A2(KEYINPUT120), .A3(new_n829), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT120), .B1(new_n791), .B2(new_n829), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT122), .B1(new_n1182), .B2(new_n246), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n792), .A2(new_n950), .B1(new_n766), .B2(new_n779), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n812), .A2(G128), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1182), .A2(KEYINPUT122), .A3(new_n246), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n770), .A2(new_n290), .B1(new_n794), .B2(new_n283), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT121), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1216), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n760), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n747), .B1(new_n835), .B2(new_n209), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n1084), .C2(new_n750), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n744), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(KEYINPUT119), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1129), .A2(new_n1130), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT119), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n744), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT123), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1233), .A2(KEYINPUT119), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1236), .B1(new_n1235), .B2(new_n744), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT123), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1232), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1136), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1235), .A2(new_n1124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1007), .A3(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(G381));
  XNOR2_X1  g1048(.A(new_n1209), .B(KEYINPUT125), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G378), .B(KEYINPUT124), .ZN(new_n1250));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n858), .A3(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(G387), .A3(G381), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G343), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1249), .A2(new_n1250), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(new_n1258), .A3(G213), .ZN(G409));
  NAND2_X1  g1059(.A1(new_n1251), .A2(G387), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G390), .B(new_n970), .C1(new_n1008), .C2(new_n991), .ZN(new_n1261));
  XOR2_X1   g1061(.A(G393), .B(G396), .Z(new_n1262));
  AND3_X1   g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1140), .B1(new_n1142), .B2(new_n1141), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1149), .B1(new_n1267), .B2(new_n1244), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1147), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1143), .A2(KEYINPUT118), .A3(new_n1149), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT57), .B1(new_n1271), .B2(new_n1170), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1174), .A2(new_n690), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1208), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1007), .B(new_n1170), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1176), .A3(new_n1202), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1250), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1257), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1257), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1245), .B1(new_n1136), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1235), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n690), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1243), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(G384), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1243), .A2(new_n858), .A3(new_n1285), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1281), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1243), .A2(new_n858), .A3(new_n1285), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n858), .B1(new_n1243), .B2(new_n1285), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1281), .B(new_n1290), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1280), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1278), .A2(new_n1279), .A3(new_n1289), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1257), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1289), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1266), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT63), .B1(new_n1302), .B2(new_n1289), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1265), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1290), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(G2897), .A3(new_n1257), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1294), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1311), .B(new_n1298), .C1(new_n1302), .C2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1306), .A2(new_n1317), .ZN(G405));
  INV_X1    g1118(.A(new_n1250), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1274), .B1(new_n1209), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1288), .A3(new_n1287), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1274), .B(new_n1289), .C1(new_n1209), .C2(new_n1319), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1321), .A2(new_n1265), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1265), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(G402));
endmodule


