//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n189), .B(new_n190), .C1(new_n192), .C2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G146), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT0), .A4(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n201), .B2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n201), .C2(G107), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G104), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n206), .A3(G104), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n206), .A3(KEYINPUT76), .A4(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n200), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n199), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n215), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n207), .B1(new_n202), .B2(new_n203), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n215), .A2(new_n200), .A3(new_n205), .A4(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(G128), .B(new_n226), .C1(new_n192), .C2(new_n194), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n196), .B(new_n197), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n201), .A2(G107), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n231), .B2(new_n207), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n218), .A2(new_n224), .B1(new_n225), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G137), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n238), .B2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n236), .A2(G134), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n241), .ZN(new_n246));
  AOI211_X1 g060(.A(G131), .B(new_n240), .C1(new_n243), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n246), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n237), .A2(new_n239), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n235), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n245), .B1(new_n244), .B2(new_n241), .ZN(new_n253));
  AOI211_X1 g067(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n236), .C2(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n249), .A2(new_n248), .A3(new_n250), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT77), .B1(new_n233), .B2(new_n225), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n223), .A2(new_n230), .A3(new_n232), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT10), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n234), .A2(new_n259), .A3(new_n260), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n252), .A2(new_n265), .A3(new_n258), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n223), .A2(new_n232), .B1(new_n229), .B2(new_n227), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n256), .A2(new_n257), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n261), .B2(new_n267), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n266), .A2(new_n268), .B1(new_n270), .B2(KEYINPUT12), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n264), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n199), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n217), .B(G101), .C1(new_n219), .C2(new_n220), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n223), .A2(KEYINPUT4), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n216), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n233), .A2(new_n225), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n263), .A2(new_n281), .A3(new_n260), .A4(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n259), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n264), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n275), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n264), .A2(new_n271), .A3(new_n276), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT79), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n187), .B(new_n188), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n264), .A2(new_n271), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n275), .B(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n285), .A2(new_n264), .A3(new_n276), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n293), .B1(new_n298), .B2(new_n187), .ZN(new_n299));
  INV_X1    g113(.A(new_n297), .ZN(new_n300));
  INV_X1    g114(.A(new_n295), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n264), .B2(new_n271), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n188), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT78), .A3(G469), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n191), .A2(G128), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n228), .A2(G143), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G134), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n238), .ZN(new_n310));
  XNOR2_X1  g124(.A(G116), .B(G122), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n309), .A2(new_n310), .B1(new_n206), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G122), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(G122), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n313), .B(new_n315), .C1(new_n316), .C2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g131(.A(G122), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT14), .B1(new_n318), .B2(G116), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(G116), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT86), .B1(new_n315), .B2(KEYINPUT14), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n317), .B(G107), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n311), .A2(new_n206), .ZN(new_n325));
  OAI21_X1  g139(.A(G107), .B1(new_n316), .B2(new_n320), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT13), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n228), .B2(G143), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n307), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n306), .A2(new_n328), .ZN(new_n331));
  OAI21_X1  g145(.A(G134), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n332), .A3(new_n310), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT68), .B(G217), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT9), .B(G234), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n334), .A2(new_n335), .A3(G953), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n324), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n324), .A2(new_n333), .ZN(new_n340));
  INV_X1    g154(.A(new_n336), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n324), .A2(new_n333), .A3(KEYINPUT87), .A4(new_n336), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT89), .B1(new_n344), .B2(new_n188), .ZN(new_n345));
  INV_X1    g159(.A(G478), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT15), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(KEYINPUT88), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(KEYINPUT88), .B2(new_n347), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n188), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n351), .B1(new_n354), .B2(new_n350), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(KEYINPUT90), .A2(G952), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT90), .A2(G952), .ZN(new_n358));
  AOI21_X1  g172(.A(G953), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G234), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT21), .B(G898), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT91), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI211_X1 g180(.A(new_n188), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  XOR2_X1   g183(.A(G113), .B(G122), .Z(new_n370));
  XOR2_X1   g184(.A(KEYINPUT84), .B(G104), .Z(new_n371));
  XOR2_X1   g185(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g186(.A(KEYINPUT16), .ZN(new_n373));
  INV_X1    g187(.A(G140), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(G125), .ZN(new_n376));
  INV_X1    g190(.A(G125), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(G146), .B(new_n375), .C1(new_n379), .C2(new_n373), .ZN(new_n380));
  NOR2_X1   g194(.A1(G237), .A2(G953), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n381), .A2(G143), .A3(G214), .ZN(new_n382));
  AOI21_X1  g196(.A(G143), .B1(new_n381), .B2(G214), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n191), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(G143), .A3(G214), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n248), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n379), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT83), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT19), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(KEYINPUT19), .B2(new_n379), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n380), .B(new_n389), .C1(new_n395), .C2(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n393), .A3(G146), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n193), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n386), .A2(new_n387), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT18), .B(G131), .C1(new_n382), .C2(new_n383), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n372), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT17), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n384), .A2(new_n388), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n375), .B1(new_n379), .B2(new_n373), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n193), .ZN(new_n408));
  OAI211_X1 g222(.A(KEYINPUT17), .B(G131), .C1(new_n382), .C2(new_n383), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n380), .A4(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n410), .A2(new_n403), .A3(new_n372), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n369), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT20), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n369), .C1(new_n404), .C2(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n372), .B1(new_n410), .B2(new_n403), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n410), .A2(new_n403), .ZN(new_n420));
  INV_X1    g234(.A(new_n372), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT85), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n419), .B1(new_n423), .B2(new_n411), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G475), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n356), .A2(new_n368), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n430));
  INV_X1    g244(.A(G119), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n314), .A2(G119), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n432), .A2(KEYINPUT5), .ZN(new_n436));
  INV_X1    g250(.A(G113), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT2), .B(G113), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n435), .A2(new_n438), .B1(new_n440), .B2(new_n434), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n223), .A3(new_n232), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n280), .A2(new_n216), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n434), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n433), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n439), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n279), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n442), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT80), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(new_n442), .C1(new_n443), .C2(new_n448), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n224), .A2(new_n447), .A3(new_n279), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n452), .B1(new_n457), .B2(new_n442), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n430), .B(new_n454), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n449), .A2(new_n453), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n455), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n377), .B1(new_n195), .B2(new_n198), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G125), .B1(new_n227), .B2(new_n229), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n467), .B(new_n469), .Z(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G210), .B1(G237), .B2(G902), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n452), .B(KEYINPUT8), .ZN(new_n475));
  INV_X1    g289(.A(new_n442), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n441), .B1(new_n223), .B2(new_n232), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n463), .A2(new_n465), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT7), .B1(new_n468), .B2(G953), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n455), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n474), .B(new_n188), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n188), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT82), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n472), .A2(new_n473), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n473), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n484), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n470), .B1(new_n459), .B2(new_n461), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n429), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G221), .B1(new_n335), .B2(G902), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n305), .A2(new_n427), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n252), .A2(new_n278), .A3(new_n258), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n244), .A2(new_n239), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G131), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n230), .A2(new_n257), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n500));
  INV_X1    g314(.A(new_n498), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n199), .B1(new_n256), .B2(new_n257), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n447), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n447), .B(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n495), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(G101), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n381), .A2(G210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n504), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT31), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT31), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n504), .A2(new_n516), .A3(new_n507), .A4(new_n513), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n447), .B1(new_n501), .B2(new_n502), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n507), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n512), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n515), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(G472), .A2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n507), .A2(new_n518), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n507), .A2(new_n520), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n513), .B(new_n528), .C1(new_n529), .C2(new_n518), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n504), .A2(new_n507), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n512), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n495), .A2(new_n498), .A3(new_n506), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n506), .B1(new_n495), .B2(new_n498), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n512), .A2(new_n533), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n528), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n188), .ZN(new_n540));
  OAI21_X1  g354(.A(G472), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n523), .A2(KEYINPUT32), .A3(new_n524), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n334), .B1(G234), .B2(new_n188), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT69), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT72), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT22), .B(G137), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OR3_X1    g364(.A1(new_n431), .A2(KEYINPUT70), .A3(G128), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT70), .B1(new_n431), .B2(G128), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(new_n552), .C1(G119), .C2(new_n228), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT24), .B(G110), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT71), .B1(new_n431), .B2(G128), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n556), .A2(KEYINPUT23), .B1(new_n431), .B2(G128), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(KEYINPUT23), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n555), .B1(new_n558), .B2(G110), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n380), .A3(new_n398), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n408), .A2(new_n380), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(G110), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(new_n562), .C1(new_n554), .C2(new_n553), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n550), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n563), .A3(new_n550), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT25), .B1(new_n567), .B2(new_n188), .ZN(new_n568));
  INV_X1    g382(.A(new_n566), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT25), .B(new_n188), .C1(new_n569), .C2(new_n564), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n546), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n544), .A2(G902), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n573), .B(KEYINPUT73), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n543), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n494), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT92), .B(G101), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G3));
  NAND2_X1  g395(.A1(new_n523), .A2(new_n188), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n582), .A2(G472), .B1(new_n524), .B2(new_n523), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n305), .A2(new_n577), .A3(new_n493), .A4(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n368), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n346), .A2(G902), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n336), .B1(new_n324), .B2(new_n333), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n324), .A2(new_n333), .A3(new_n336), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(KEYINPUT93), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n337), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n339), .A2(new_n342), .A3(new_n587), .A4(new_n343), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n586), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT94), .B(G478), .Z(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n344), .B2(new_n188), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n416), .A2(new_n425), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n492), .A2(new_n585), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n584), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT34), .B(G104), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  NOR2_X1   g418(.A1(new_n355), .A2(new_n426), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n492), .A2(new_n585), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n584), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G107), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  NAND2_X1  g424(.A1(new_n560), .A2(new_n563), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n574), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n572), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n572), .A2(KEYINPUT96), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n583), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n494), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT37), .B(G110), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G12));
  INV_X1    g438(.A(G900), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n363), .B1(new_n625), .B2(new_n367), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n355), .A2(new_n426), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n305), .A2(new_n492), .A3(new_n493), .A4(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT29), .B1(new_n531), .B2(new_n512), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n540), .B1(new_n530), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G472), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n542), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT32), .B1(new_n523), .B2(new_n524), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n619), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n228), .ZN(G30));
  NAND2_X1  g450(.A1(new_n487), .A2(new_n491), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n487), .A2(KEYINPUT38), .A3(new_n491), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n495), .A2(new_n498), .ZN(new_n642));
  INV_X1    g456(.A(new_n506), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n507), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n188), .B1(new_n645), .B2(new_n513), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n512), .B1(new_n504), .B2(new_n507), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n527), .A2(new_n542), .A3(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n413), .A2(new_n415), .B1(new_n424), .B2(G475), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n355), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n619), .A2(new_n429), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n641), .A2(new_n649), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n305), .A2(new_n493), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n626), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(KEYINPUT40), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n653), .A2(new_n654), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n655), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  INV_X1    g480(.A(new_n626), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n600), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n324), .A2(new_n333), .A3(KEYINPUT93), .A4(new_n336), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n342), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n337), .A2(new_n591), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT33), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n594), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n598), .B1(new_n673), .B2(new_n586), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n650), .A2(new_n674), .A3(KEYINPUT99), .A4(new_n626), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n305), .A2(new_n676), .A3(new_n492), .A4(new_n493), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(new_n634), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n287), .A2(new_n288), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n291), .B1(new_n681), .B2(new_n290), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n680), .B(G469), .C1(new_n682), .C2(G902), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n276), .B1(new_n285), .B2(new_n264), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n290), .B1(new_n684), .B2(KEYINPUT79), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n277), .A2(new_n288), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT100), .B1(new_n687), .B2(new_n187), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n493), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n687), .B2(new_n187), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n689), .A2(new_n577), .A3(new_n543), .A4(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(new_n692), .B2(new_n601), .ZN(new_n693));
  INV_X1    g507(.A(new_n601), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n523), .A2(KEYINPUT32), .A3(new_n524), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n519), .B1(new_n645), .B2(KEYINPUT28), .ZN(new_n696));
  AOI21_X1  g510(.A(G902), .B1(new_n696), .B2(new_n538), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n629), .A2(new_n530), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n631), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n576), .B1(new_n700), .B2(new_n527), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n292), .A2(new_n493), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n683), .B2(new_n688), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n694), .A2(new_n701), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n693), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  AND3_X1   g522(.A1(new_n492), .A2(new_n585), .A3(new_n605), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n701), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AOI22_X1  g525(.A1(new_n700), .A2(new_n527), .B1(new_n617), .B2(new_n618), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n703), .A3(new_n427), .A4(new_n492), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  AND3_X1   g528(.A1(new_n492), .A2(new_n585), .A3(new_n651), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n631), .B1(new_n523), .B2(new_n188), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n514), .A2(KEYINPUT31), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n513), .B1(new_n537), .B2(new_n528), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT102), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n515), .B(new_n720), .C1(new_n696), .C2(new_n513), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n517), .A3(new_n721), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n576), .B(new_n716), .C1(new_n722), .C2(new_n524), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n703), .A2(new_n715), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NAND2_X1  g539(.A1(new_n685), .A2(new_n686), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n188), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n680), .B1(new_n727), .B2(G469), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n687), .A2(KEYINPUT100), .A3(new_n187), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n492), .B(new_n691), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n722), .A2(new_n524), .ZN(new_n731));
  INV_X1    g545(.A(new_n716), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n676), .A3(new_n732), .A4(new_n619), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n377), .ZN(G27));
  NOR2_X1   g549(.A1(new_n690), .A2(new_n429), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n487), .A2(new_n491), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n303), .A2(G469), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n292), .A2(new_n738), .ZN(new_n739));
  AND4_X1   g553(.A1(KEYINPUT42), .A2(new_n737), .A3(new_n676), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n700), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n740), .A2(new_n741), .A3(new_n577), .A4(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n541), .B(new_n542), .C1(KEYINPUT103), .C2(new_n633), .ZN(new_n746));
  INV_X1    g560(.A(new_n743), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n577), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n737), .A2(new_n676), .A3(new_n739), .A4(KEYINPUT42), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT104), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT105), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n487), .A2(new_n491), .A3(new_n736), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n292), .B2(new_n738), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n701), .A2(new_n676), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n752), .B1(new_n751), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT106), .B(G131), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G33));
  NAND3_X1  g576(.A1(new_n701), .A2(new_n627), .A3(new_n754), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  AND2_X1   g578(.A1(new_n617), .A2(new_n618), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT43), .B1(new_n426), .B2(new_n674), .ZN(new_n766));
  INV_X1    g580(.A(new_n674), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n650), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n765), .A2(new_n583), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n772));
  AOI211_X1 g586(.A(G469), .B(G902), .C1(new_n685), .C2(new_n686), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n300), .B2(new_n302), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n296), .A2(KEYINPUT45), .A3(new_n297), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(G469), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(new_n493), .A3(new_n657), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n487), .A2(new_n428), .A3(new_n491), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT107), .Z(new_n787));
  NAND4_X1  g601(.A1(new_n772), .A2(new_n784), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  AND2_X1   g603(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n790));
  NOR2_X1   g604(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n783), .B2(new_n493), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n690), .B(new_n790), .C1(new_n781), .C2(new_n782), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n676), .A2(new_n576), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n786), .A3(new_n543), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  OR2_X1    g613(.A1(G952), .A2(G953), .ZN(new_n800));
  XNOR2_X1  g614(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n428), .B1(new_n639), .B2(new_n640), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n703), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n770), .A2(new_n362), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n723), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n801), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n649), .A2(new_n576), .A3(new_n362), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n773), .B1(new_n683), .B2(new_n688), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n767), .A2(new_n426), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n737), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n716), .B1(new_n722), .B2(new_n524), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(new_n577), .A3(new_n804), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(KEYINPUT50), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n703), .A3(new_n814), .A4(new_n802), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n731), .A2(new_n732), .A3(new_n619), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n737), .A3(new_n808), .A4(new_n804), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n806), .A2(new_n810), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT116), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n810), .A2(new_n817), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n815), .A4(new_n806), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n689), .A2(KEYINPUT114), .A3(new_n292), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n690), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n793), .A2(new_n794), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n787), .A2(new_n812), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n819), .A2(new_n822), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n819), .A2(new_n822), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n808), .A2(new_n737), .A3(new_n804), .ZN(new_n835));
  INV_X1    g649(.A(new_n748), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT48), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n807), .A2(new_n600), .A3(new_n737), .A4(new_n808), .ZN(new_n839));
  INV_X1    g653(.A(new_n730), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n812), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n359), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n827), .A2(new_n828), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n820), .A3(new_n815), .A4(new_n806), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n823), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n834), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n834), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n713), .A2(new_n710), .A3(new_n724), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n584), .B1(new_n601), .B2(new_n606), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n579), .A3(new_n621), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n786), .A2(new_n356), .A3(new_n426), .A4(new_n626), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n712), .A2(new_n854), .A3(new_n656), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n754), .A2(new_n619), .A3(new_n676), .A4(new_n811), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n855), .A2(new_n763), .A3(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n706), .A2(new_n851), .A3(new_n853), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n759), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n745), .A2(new_n750), .B1(new_n756), .B2(new_n755), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n752), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n730), .A2(new_n733), .B1(new_n628), .B2(new_n634), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n615), .A2(new_n690), .A3(new_n626), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n739), .A2(new_n492), .A3(new_n651), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n649), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n677), .A2(new_n634), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n862), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n862), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n858), .A2(new_n859), .A3(new_n861), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n862), .A2(KEYINPUT112), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT112), .ZN(new_n875));
  OAI221_X1 g689(.A(new_n875), .B1(new_n628), .B2(new_n634), .C1(new_n730), .C2(new_n733), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n864), .A2(new_n865), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n867), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n874), .A2(new_n876), .A3(new_n678), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n869), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n760), .A2(new_n873), .A3(new_n858), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(KEYINPUT54), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n873), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n691), .B1(new_n728), .B2(new_n729), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n578), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n543), .A2(new_n427), .A3(new_n619), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n887), .A2(new_n709), .B1(new_n840), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n706), .A2(new_n889), .A3(new_n724), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n885), .B1(new_n890), .B2(new_n860), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n751), .A2(new_n757), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT113), .A3(new_n706), .A4(new_n851), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n853), .A2(new_n857), .A3(KEYINPUT53), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n869), .B2(new_n879), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n883), .A2(new_n884), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n882), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n800), .B1(new_n850), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n577), .A2(new_n736), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT109), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n650), .B(new_n767), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT110), .Z(new_n905));
  NOR3_X1   g719(.A1(new_n905), .A2(new_n649), .A3(new_n641), .ZN(new_n906));
  INV_X1    g720(.A(new_n808), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(KEYINPUT49), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(KEYINPUT49), .B2(new_n907), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT111), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n900), .A2(new_n910), .ZN(G75));
  NOR2_X1   g725(.A1(new_n273), .A2(G952), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT120), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n462), .B(KEYINPUT119), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n470), .B(KEYINPUT55), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n915), .B(new_n916), .Z(new_n917));
  AOI22_X1  g731(.A1(new_n873), .A2(new_n871), .B1(new_n894), .B2(new_n896), .ZN(new_n918));
  INV_X1    g732(.A(G210), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n188), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n920), .B2(KEYINPUT56), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  INV_X1    g736(.A(new_n917), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n883), .A2(new_n897), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G902), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n923), .C1(new_n925), .C2(new_n919), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n914), .B1(new_n921), .B2(new_n926), .ZN(G51));
  XOR2_X1   g741(.A(new_n778), .B(KEYINPUT57), .Z(new_n928));
  AND3_X1   g742(.A1(new_n883), .A2(new_n884), .A3(new_n897), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n884), .B1(new_n883), .B2(new_n897), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n726), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n777), .B(KEYINPUT121), .Z(new_n933));
  NAND3_X1  g747(.A1(new_n924), .A2(G902), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n912), .B1(new_n932), .B2(new_n934), .ZN(G54));
  NOR2_X1   g749(.A1(new_n404), .A2(new_n411), .ZN(new_n936));
  NAND2_X1  g750(.A1(KEYINPUT58), .A2(G475), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n925), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n912), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n925), .A2(new_n936), .A3(new_n937), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(G60));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n673), .B1(new_n899), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n673), .A2(new_n945), .ZN(new_n947));
  INV_X1    g761(.A(new_n930), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n898), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n946), .A2(new_n949), .A3(new_n914), .ZN(G63));
  INV_X1    g764(.A(new_n567), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT122), .Z(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n951), .B1(new_n918), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n883), .B2(new_n897), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n914), .B1(new_n957), .B2(new_n613), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n957), .B2(new_n613), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n956), .B(new_n958), .C1(new_n960), .C2(KEYINPUT61), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n851), .A2(new_n853), .A3(new_n857), .A4(new_n706), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n962), .A2(new_n758), .A3(new_n759), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT53), .B1(new_n963), .B2(new_n870), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n853), .A2(new_n857), .A3(KEYINPUT53), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n880), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n891), .B2(new_n893), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n613), .B(new_n954), .C1(new_n964), .C2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT61), .B1(new_n968), .B2(KEYINPUT123), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n956), .A2(new_n913), .A3(new_n968), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n961), .A2(new_n971), .ZN(G66));
  AOI21_X1  g786(.A(new_n273), .B1(new_n365), .B2(G224), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n851), .A2(new_n853), .A3(new_n706), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n273), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n915), .B1(G898), .B2(new_n273), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT124), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  NAND2_X1  g792(.A1(G227), .A2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n499), .A2(new_n503), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(new_n395), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n874), .A2(new_n678), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n876), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n798), .A2(new_n788), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n784), .A2(new_n492), .A3(new_n651), .A4(new_n836), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n986), .A2(new_n763), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n760), .A2(new_n984), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n273), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n625), .A2(G953), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT126), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n982), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n984), .A2(new_n994), .A3(new_n664), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n605), .A2(new_n600), .ZN(new_n996));
  OR4_X1    g810(.A1(new_n578), .A2(new_n658), .A3(new_n786), .A4(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n985), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n664), .A2(new_n983), .A3(new_n876), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n995), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n995), .A2(new_n998), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n980), .B(new_n993), .C1(new_n1005), .C2(new_n982), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n989), .A2(new_n992), .ZN(new_n1007));
  INV_X1    g821(.A(new_n982), .ZN(new_n1008));
  OAI211_X1 g822(.A(G953), .B(new_n979), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n988), .B2(new_n974), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1013), .A2(new_n507), .A3(new_n504), .A4(new_n512), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n514), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(new_n532), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n872), .A2(new_n881), .A3(new_n1012), .A4(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1014), .A2(new_n939), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1012), .B1(new_n1020), .B2(new_n974), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1019), .B1(new_n1021), .B2(new_n647), .ZN(G57));
endmodule


