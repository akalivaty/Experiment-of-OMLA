

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U323 ( .A(n412), .B(n411), .ZN(n524) );
  XNOR2_X1 U324 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U325 ( .A(n410), .B(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U326 ( .A(n371), .B(n370), .ZN(n372) );
  OR2_X1 U327 ( .A1(n428), .A2(n568), .ZN(n429) );
  XNOR2_X1 U328 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U329 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(G36GAT), .B(G190GAT), .Z(n417) );
  XOR2_X1 U331 ( .A(G99GAT), .B(G85GAT), .Z(n364) );
  XOR2_X1 U332 ( .A(n417), .B(n364), .Z(n292) );
  XOR2_X1 U333 ( .A(G50GAT), .B(G162GAT), .Z(n336) );
  XOR2_X1 U334 ( .A(G134GAT), .B(KEYINPUT75), .Z(n323) );
  XNOR2_X1 U335 ( .A(n336), .B(n323), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U337 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U338 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n350) );
  XOR2_X1 U340 ( .A(G92GAT), .B(n350), .Z(n296) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U343 ( .A(n298), .B(n297), .Z(n306) );
  XOR2_X1 U344 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n300) );
  XNOR2_X1 U345 ( .A(G218GAT), .B(KEYINPUT67), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U347 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n302) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n554) );
  XOR2_X1 U352 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n308) );
  XNOR2_X1 U353 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(G141GAT), .B(n309), .Z(n335) );
  XOR2_X1 U356 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n311) );
  XNOR2_X1 U357 ( .A(G1GAT), .B(KEYINPUT91), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U359 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n313) );
  XNOR2_X1 U360 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U362 ( .A(n315), .B(n314), .Z(n329) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G127GAT), .Z(n317) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n433) );
  XOR2_X1 U366 ( .A(n433), .B(KEYINPUT89), .Z(n319) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n327) );
  XOR2_X1 U369 ( .A(G57GAT), .B(G155GAT), .Z(n321) );
  XNOR2_X1 U370 ( .A(G148GAT), .B(G162GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(n322), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U377 ( .A(n335), .B(n330), .Z(n511) );
  XNOR2_X1 U378 ( .A(G211GAT), .B(KEYINPUT84), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n331), .B(KEYINPUT21), .ZN(n332) );
  XOR2_X1 U380 ( .A(n332), .B(KEYINPUT85), .Z(n334) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U382 ( .A(n334), .B(n333), .ZN(n423) );
  XNOR2_X1 U383 ( .A(n423), .B(n335), .ZN(n347) );
  XOR2_X1 U384 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n338) );
  XOR2_X1 U385 ( .A(G22GAT), .B(G155GAT), .Z(n390) );
  XNOR2_X1 U386 ( .A(n336), .B(n390), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U388 ( .A(n339), .B(KEYINPUT23), .Z(n345) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n340), .B(G148GAT), .ZN(n371) );
  XOR2_X1 U391 ( .A(KEYINPUT24), .B(n371), .Z(n342) );
  NAND2_X1 U392 ( .A1(G228GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n343), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n460) );
  NAND2_X1 U397 ( .A1(n511), .A2(n460), .ZN(n428) );
  INV_X1 U398 ( .A(KEYINPUT54), .ZN(n427) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G197GAT), .Z(n349) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G22GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n363) );
  XOR2_X1 U402 ( .A(G15GAT), .B(G1GAT), .Z(n398) );
  XOR2_X1 U403 ( .A(n398), .B(G36GAT), .Z(n352) );
  XNOR2_X1 U404 ( .A(n350), .B(G50GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U406 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n354) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U409 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U410 ( .A(KEYINPUT29), .B(G8GAT), .Z(n358) );
  XNOR2_X1 U411 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n359), .B(KEYINPUT70), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n543) );
  INV_X1 U416 ( .A(n543), .ZN(n572) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(n364), .ZN(n365) );
  XOR2_X1 U418 ( .A(n365), .B(KEYINPUT31), .Z(n380) );
  XOR2_X1 U419 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n367) );
  XNOR2_X1 U420 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n373) );
  NAND2_X1 U422 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  INV_X1 U423 ( .A(KEYINPUT73), .ZN(n368) );
  XOR2_X1 U424 ( .A(n373), .B(n372), .Z(n378) );
  XNOR2_X1 U425 ( .A(G71GAT), .B(G57GAT), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n374), .B(KEYINPUT13), .ZN(n387) );
  XOR2_X1 U427 ( .A(G64GAT), .B(G92GAT), .Z(n376) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G204GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n422) );
  XNOR2_X1 U430 ( .A(n387), .B(n422), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n576) );
  XOR2_X1 U433 ( .A(KEYINPUT41), .B(n576), .Z(n545) );
  NOR2_X1 U434 ( .A1(n572), .A2(n545), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n381), .B(KEYINPUT112), .ZN(n383) );
  INV_X1 U436 ( .A(KEYINPUT46), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n403) );
  XOR2_X1 U438 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n389) );
  XOR2_X1 U439 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n385) );
  XNOR2_X1 U440 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n394) );
  XOR2_X1 U444 ( .A(G8GAT), .B(G183GAT), .Z(n420) );
  XOR2_X1 U445 ( .A(n420), .B(n390), .Z(n392) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U448 ( .A(n394), .B(n393), .Z(n400) );
  XOR2_X1 U449 ( .A(G64GAT), .B(G78GAT), .Z(n396) );
  XNOR2_X1 U450 ( .A(G127GAT), .B(G211GAT), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U453 ( .A(n400), .B(n399), .Z(n581) );
  XNOR2_X1 U454 ( .A(n581), .B(KEYINPUT111), .ZN(n564) );
  INV_X1 U455 ( .A(n554), .ZN(n401) );
  NOR2_X1 U456 ( .A1(n564), .A2(n401), .ZN(n402) );
  NAND2_X1 U457 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n404), .B(KEYINPUT47), .ZN(n409) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(n554), .ZN(n584) );
  NOR2_X1 U460 ( .A1(n584), .A2(n581), .ZN(n405) );
  XNOR2_X1 U461 ( .A(KEYINPUT45), .B(n405), .ZN(n406) );
  NAND2_X1 U462 ( .A1(n406), .A2(n576), .ZN(n407) );
  NOR2_X1 U463 ( .A1(n543), .A2(n407), .ZN(n408) );
  NOR2_X1 U464 ( .A1(n409), .A2(n408), .ZN(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n410) );
  XNOR2_X1 U466 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n413), .B(KEYINPUT82), .ZN(n414) );
  XOR2_X1 U468 ( .A(n414), .B(KEYINPUT81), .Z(n416) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n415) );
  XOR2_X1 U470 ( .A(n416), .B(n415), .Z(n444) );
  XNOR2_X1 U471 ( .A(n417), .B(n444), .ZN(n419) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U474 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U476 ( .A(n425), .B(n424), .Z(n488) );
  INV_X1 U477 ( .A(n488), .ZN(n514) );
  NOR2_X1 U478 ( .A1(n524), .A2(n514), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n568) );
  XNOR2_X1 U480 ( .A(n429), .B(KEYINPUT120), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n430), .B(KEYINPUT55), .ZN(n446) );
  XOR2_X1 U482 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U483 ( .A(G176GAT), .B(G71GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n443) );
  XOR2_X1 U485 ( .A(G99GAT), .B(n433), .Z(n435) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G190GAT), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U488 ( .A(n436), .B(G134GAT), .Z(n441) );
  XOR2_X1 U489 ( .A(G183GAT), .B(KEYINPUT79), .Z(n438) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U495 ( .A(n445), .B(n444), .Z(n516) );
  INV_X1 U496 ( .A(n516), .ZN(n526) );
  NAND2_X1 U497 ( .A1(n446), .A2(n526), .ZN(n563) );
  NOR2_X1 U498 ( .A1(n554), .A2(n563), .ZN(n450) );
  XNOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n448) );
  INV_X1 U500 ( .A(G190GAT), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n452) );
  XNOR2_X1 U502 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n469) );
  AND2_X1 U504 ( .A1(n543), .A2(n576), .ZN(n482) );
  NAND2_X1 U505 ( .A1(n526), .A2(n488), .ZN(n453) );
  NAND2_X1 U506 ( .A1(n460), .A2(n453), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT25), .B(n454), .Z(n458) );
  NOR2_X1 U508 ( .A1(n460), .A2(n526), .ZN(n456) );
  XNOR2_X1 U509 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n570) );
  XNOR2_X1 U511 ( .A(n488), .B(KEYINPUT27), .ZN(n462) );
  NAND2_X1 U512 ( .A1(n570), .A2(n462), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n511), .A2(n459), .ZN(n465) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT68), .ZN(n461) );
  XOR2_X1 U516 ( .A(n461), .B(KEYINPUT28), .Z(n494) );
  INV_X1 U517 ( .A(n494), .ZN(n527) );
  INV_X1 U518 ( .A(n511), .ZN(n569) );
  NAND2_X1 U519 ( .A1(n462), .A2(n569), .ZN(n523) );
  NOR2_X1 U520 ( .A1(n526), .A2(n523), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n527), .A2(n463), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n478) );
  INV_X1 U523 ( .A(n581), .ZN(n550) );
  NAND2_X1 U524 ( .A1(n554), .A2(n550), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n466), .Z(n467) );
  AND2_X1 U526 ( .A1(n478), .A2(n467), .ZN(n499) );
  NAND2_X1 U527 ( .A1(n482), .A2(n499), .ZN(n474) );
  NOR2_X1 U528 ( .A1(n511), .A2(n474), .ZN(n468) );
  XOR2_X1 U529 ( .A(n469), .B(n468), .Z(G1324GAT) );
  NOR2_X1 U530 ( .A1(n514), .A2(n474), .ZN(n471) );
  XNOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U533 ( .A1(n516), .A2(n474), .ZN(n473) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n473), .B(n472), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n527), .A2(n474), .ZN(n476) );
  XNOR2_X1 U537 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n477), .ZN(G1327GAT) );
  NAND2_X1 U540 ( .A1(n581), .A2(n478), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n584), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT99), .B(KEYINPUT37), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n510) );
  NAND2_X1 U544 ( .A1(n482), .A2(n510), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n483), .Z(n495) );
  NAND2_X1 U546 ( .A1(n495), .A2(n569), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n485) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT98), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n495), .A2(n488), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n491) );
  NAND2_X1 U555 ( .A1(n495), .A2(n526), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1330GAT) );
  XOR2_X1 U558 ( .A(G50GAT), .B(KEYINPUT103), .Z(n497) );
  NAND2_X1 U559 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(n545), .B(KEYINPUT105), .Z(n558) );
  NOR2_X1 U562 ( .A1(n543), .A2(n558), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(KEYINPUT106), .ZN(n509) );
  NAND2_X1 U564 ( .A1(n499), .A2(n509), .ZN(n505) );
  NOR2_X1 U565 ( .A1(n511), .A2(n505), .ZN(n501) );
  XNOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n505), .ZN(n503) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n516), .A2(n505), .ZN(n504) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n527), .A2(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  NAND2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n519) );
  NOR2_X1 U578 ( .A1(n511), .A2(n519), .ZN(n512) );
  XOR2_X1 U579 ( .A(n512), .B(KEYINPUT108), .Z(n513) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n519), .ZN(n515) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n519), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n527), .A2(n519), .ZN(n521) );
  XNOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n522), .Z(G1339GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT114), .B(n525), .ZN(n542) );
  AND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n542), .A2(n528), .ZN(n537) );
  INV_X1 U594 ( .A(n537), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n533), .A2(n543), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U597 ( .A1(n558), .A2(n537), .ZN(n531) );
  XNOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U602 ( .A1(n533), .A2(n564), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  NOR2_X1 U605 ( .A1(n537), .A2(n554), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n539) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n542), .A2(n570), .ZN(n553) );
  INV_X1 U611 ( .A(n553), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n551), .A2(n543), .ZN(n544) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  NOR2_X1 U614 ( .A1(n553), .A2(n545), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n547) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n546) );
  XNOR2_X1 U617 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n572), .A2(n563), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G169GAT), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT121), .ZN(G1348GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n563), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .Z(n567) );
  INV_X1 U632 ( .A(n563), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n583) );
  NOR2_X1 U637 ( .A1(n572), .A2(n583), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n583), .A2(n576), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

