

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U552 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X2 U553 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  NOR2_X2 U554 ( .A1(n528), .A2(n527), .ZN(G160) );
  NOR2_X1 U555 ( .A1(n957), .A2(n696), .ZN(n703) );
  XNOR2_X1 U556 ( .A(n722), .B(KEYINPUT30), .ZN(n723) );
  AND2_X1 U557 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U558 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X2 U559 ( .A(n684), .B(KEYINPUT64), .ZN(n719) );
  INV_X1 U560 ( .A(n719), .ZN(n697) );
  XNOR2_X1 U561 ( .A(n724), .B(n723), .ZN(n725) );
  INV_X1 U562 ( .A(n940), .ZN(n750) );
  INV_X1 U563 ( .A(KEYINPUT101), .ZN(n759) );
  NOR2_X1 U564 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U565 ( .A1(G651), .A2(n644), .ZN(n649) );
  INV_X1 U566 ( .A(G2104), .ZN(n519) );
  AND2_X1 U567 ( .A1(n519), .A2(G2105), .ZN(n873) );
  NAND2_X1 U568 ( .A1(n873), .A2(G125), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G2105), .A2(n519), .ZN(n529) );
  NAND2_X1 U570 ( .A1(G101), .A2(n529), .ZN(n520) );
  XOR2_X1 U571 ( .A(n520), .B(KEYINPUT23), .Z(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n528) );
  XNOR2_X2 U573 ( .A(n524), .B(n523), .ZN(n877) );
  NAND2_X1 U574 ( .A1(G137), .A2(n877), .ZN(n526) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U576 ( .A1(G113), .A2(n874), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G138), .A2(n877), .ZN(n532) );
  INV_X1 U579 ( .A(n529), .ZN(n530) );
  INV_X1 U580 ( .A(n530), .ZN(n878) );
  NAND2_X1 U581 ( .A1(G102), .A2(n878), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U583 ( .A1(G126), .A2(n873), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G114), .A2(n874), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U586 ( .A1(n536), .A2(n535), .ZN(G164) );
  XNOR2_X1 U587 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n635) );
  NAND2_X1 U589 ( .A1(G85), .A2(n635), .ZN(n538) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  INV_X1 U591 ( .A(G651), .ZN(n539) );
  NOR2_X1 U592 ( .A1(n644), .A2(n539), .ZN(n638) );
  NAND2_X1 U593 ( .A1(G72), .A2(n638), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n546) );
  NAND2_X1 U595 ( .A1(n649), .A2(G47), .ZN(n544) );
  NOR2_X1 U596 ( .A1(G543), .A2(n539), .ZN(n541) );
  XNOR2_X1 U597 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U599 ( .A(KEYINPUT66), .B(n542), .ZN(n648) );
  NAND2_X1 U600 ( .A1(G60), .A2(n648), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U602 ( .A1(n546), .A2(n545), .ZN(G290) );
  NAND2_X1 U603 ( .A1(n649), .A2(G52), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G64), .A2(n648), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G90), .A2(n635), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G77), .A2(n638), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT68), .B(n551), .Z(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n552), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n554), .A2(n553), .ZN(G171) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  NAND2_X1 U616 ( .A1(n649), .A2(G51), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G63), .A2(n648), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n557), .Z(n565) );
  NAND2_X1 U620 ( .A1(G76), .A2(n638), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n559) );
  NAND2_X1 U622 ( .A1(G89), .A2(n635), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT74), .ZN(n563) );
  XNOR2_X1 U626 ( .A(KEYINPUT5), .B(n563), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U628 ( .A(KEYINPUT7), .B(n566), .ZN(G168) );
  XNOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .ZN(n567) );
  XNOR2_X1 U630 ( .A(n567), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT10), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT70), .B(n569), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n823) );
  NAND2_X1 U635 ( .A1(n823), .A2(G567), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT71), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT11), .B(n571), .ZN(G234) );
  NAND2_X1 U638 ( .A1(n648), .A2(G56), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n572), .Z(n578) );
  NAND2_X1 U640 ( .A1(n635), .A2(G81), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G68), .A2(n638), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n649), .A2(G43), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n957) );
  INV_X1 U648 ( .A(G860), .ZN(n624) );
  OR2_X1 U649 ( .A1(n957), .A2(n624), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G54), .A2(n649), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n638), .A2(G79), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G66), .A2(n648), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n635), .A2(G92), .ZN(n583) );
  XOR2_X1 U657 ( .A(KEYINPUT72), .B(n583), .Z(n584) );
  NOR2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT15), .ZN(n942) );
  OR2_X1 U661 ( .A1(n942), .A2(G868), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G91), .A2(n635), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G78), .A2(n638), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G65), .A2(n648), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(n593), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n649), .A2(G53), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G299) );
  INV_X1 U671 ( .A(G868), .ZN(n662) );
  NOR2_X1 U672 ( .A1(G286), .A2(n662), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n624), .A2(G559), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n600), .A2(n942), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT76), .ZN(n602) );
  XNOR2_X1 U678 ( .A(KEYINPUT16), .B(n602), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n957), .ZN(n603) );
  XOR2_X1 U680 ( .A(KEYINPUT77), .B(n603), .Z(n606) );
  NAND2_X1 U681 ( .A1(G868), .A2(n942), .ZN(n604) );
  NOR2_X1 U682 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U684 ( .A(KEYINPUT78), .B(n607), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n873), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n878), .A2(G99), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G135), .A2(n877), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G111), .A2(n874), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n1001) );
  XNOR2_X1 U693 ( .A(n1001), .B(G2096), .ZN(n616) );
  INV_X1 U694 ( .A(G2100), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U696 ( .A1(n635), .A2(G93), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G67), .A2(n648), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G80), .A2(n638), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G55), .A2(n649), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n661) );
  NAND2_X1 U703 ( .A1(G559), .A2(n942), .ZN(n623) );
  XOR2_X1 U704 ( .A(n957), .B(n623), .Z(n659) );
  NAND2_X1 U705 ( .A1(n624), .A2(n659), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n625), .B(KEYINPUT79), .ZN(n626) );
  XOR2_X1 U707 ( .A(n661), .B(n626), .Z(G145) );
  NAND2_X1 U708 ( .A1(G48), .A2(n649), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n635), .A2(G86), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G61), .A2(n648), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n638), .A2(G73), .ZN(n629) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U717 ( .A1(n635), .A2(G88), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G62), .A2(n648), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G75), .A2(n638), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G50), .A2(n649), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n643), .Z(G166) );
  NAND2_X1 U725 ( .A1(G87), .A2(n644), .ZN(n646) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n649), .A2(G49), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G288) );
  XNOR2_X1 U731 ( .A(G305), .B(G166), .ZN(n658) );
  XNOR2_X1 U732 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U733 ( .A(G288), .B(KEYINPUT82), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U735 ( .A(n661), .B(n654), .Z(n656) );
  INV_X1 U736 ( .A(G299), .ZN(n946) );
  XNOR2_X1 U737 ( .A(G290), .B(n946), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U739 ( .A(n658), .B(n657), .ZN(n848) );
  XNOR2_X1 U740 ( .A(n659), .B(n848), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n660), .A2(G868), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n668), .A2(G2072), .ZN(n669) );
  XNOR2_X1 U749 ( .A(KEYINPUT84), .B(n669), .ZN(G158) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n670) );
  NOR2_X1 U751 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G108), .A2(n671), .ZN(n827) );
  NAND2_X1 U753 ( .A1(G567), .A2(n827), .ZN(n672) );
  XNOR2_X1 U754 ( .A(n672), .B(KEYINPUT85), .ZN(n677) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT22), .B(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G96), .ZN(n675) );
  OR2_X1 U758 ( .A1(G218), .A2(n675), .ZN(n828) );
  AND2_X1 U759 ( .A1(G2106), .A2(n828), .ZN(n676) );
  NOR2_X1 U760 ( .A1(n677), .A2(n676), .ZN(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n679) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n679), .A2(n678), .ZN(n826) );
  NAND2_X1 U764 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U766 ( .A(G1986), .B(KEYINPUT86), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n680), .B(G290), .ZN(n949) );
  NOR2_X2 U768 ( .A1(G164), .A2(G1384), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n681) );
  NOR2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n818) );
  NAND2_X1 U771 ( .A1(n949), .A2(n818), .ZN(n807) );
  AND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n683) );
  XOR2_X1 U773 ( .A(G2078), .B(KEYINPUT25), .Z(n917) );
  NOR2_X1 U774 ( .A1(n719), .A2(n917), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT93), .ZN(n687) );
  OR2_X1 U776 ( .A1(n697), .A2(G1961), .ZN(n686) );
  NAND2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n726) );
  NAND2_X1 U778 ( .A1(n726), .A2(G171), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n697), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U780 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n689), .B(n688), .ZN(n691) );
  XNOR2_X1 U782 ( .A(G1956), .B(KEYINPUT95), .ZN(n976) );
  NOR2_X1 U783 ( .A1(n697), .A2(n976), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n706) );
  NOR2_X1 U785 ( .A1(n946), .A2(n706), .ZN(n692) );
  XOR2_X1 U786 ( .A(n692), .B(KEYINPUT28), .Z(n710) );
  NAND2_X1 U787 ( .A1(n719), .A2(G1341), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n697), .A2(G1996), .ZN(n693) );
  XNOR2_X1 U789 ( .A(n693), .B(KEYINPUT26), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n942), .A2(n703), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n697), .A2(G2067), .ZN(n698) );
  XNOR2_X1 U793 ( .A(n698), .B(KEYINPUT96), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n719), .A2(G1348), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n705) );
  OR2_X1 U797 ( .A1(n942), .A2(n703), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U799 ( .A1(n946), .A2(n706), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U802 ( .A(n711), .B(KEYINPUT29), .Z(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n738) );
  INV_X1 U804 ( .A(G8), .ZN(n718) );
  NOR2_X1 U805 ( .A1(n719), .A2(G2090), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n719), .A2(G8), .ZN(n771) );
  NOR2_X1 U807 ( .A1(G1971), .A2(n771), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n716), .A2(G303), .ZN(n717) );
  OR2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n732) );
  AND2_X1 U811 ( .A1(n738), .A2(n732), .ZN(n731) );
  INV_X1 U812 ( .A(KEYINPUT31), .ZN(n730) );
  NOR2_X1 U813 ( .A1(n719), .A2(G2084), .ZN(n741) );
  NOR2_X1 U814 ( .A1(n771), .A2(G1966), .ZN(n720) );
  XNOR2_X1 U815 ( .A(n720), .B(KEYINPUT92), .ZN(n740) );
  NOR2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n721), .A2(G8), .ZN(n724) );
  XOR2_X1 U818 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n722) );
  NOR2_X1 U819 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U820 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n730), .B(n729), .ZN(n739) );
  NAND2_X1 U823 ( .A1(n731), .A2(n739), .ZN(n736) );
  INV_X1 U824 ( .A(n732), .ZN(n734) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n733) );
  OR2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U828 ( .A(n737), .B(KEYINPUT32), .ZN(n748) );
  AND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n745) );
  INV_X1 U830 ( .A(n740), .ZN(n743) );
  NAND2_X1 U831 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U834 ( .A(n746), .B(KEYINPUT99), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n764) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n754), .A2(n749), .ZN(n955) );
  NAND2_X1 U839 ( .A1(n764), .A2(n955), .ZN(n752) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n940) );
  NOR2_X1 U841 ( .A1(n771), .A2(n750), .ZN(n751) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n753), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  XNOR2_X1 U844 ( .A(KEYINPUT100), .B(n755), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n756), .A2(n771), .ZN(n757) );
  NOR2_X2 U846 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U847 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n936) );
  NAND2_X1 U849 ( .A1(n761), .A2(n936), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n765), .A2(n771), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT102), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U857 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n805) );
  XNOR2_X1 U860 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G128), .A2(n873), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G116), .A2(n874), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n777), .B(n776), .ZN(n784) );
  NAND2_X1 U865 ( .A1(n877), .A2(G140), .ZN(n778) );
  XOR2_X1 U866 ( .A(KEYINPUT87), .B(n778), .Z(n780) );
  NAND2_X1 U867 ( .A1(n878), .A2(G104), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n782) );
  XOR2_X1 U869 ( .A(KEYINPUT88), .B(KEYINPUT34), .Z(n781) );
  XOR2_X1 U870 ( .A(n782), .B(n781), .Z(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U872 ( .A(KEYINPUT36), .B(n785), .ZN(n893) );
  XNOR2_X1 U873 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NOR2_X1 U874 ( .A1(n893), .A2(n815), .ZN(n1017) );
  NAND2_X1 U875 ( .A1(n818), .A2(n1017), .ZN(n813) );
  NAND2_X1 U876 ( .A1(G131), .A2(n877), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G119), .A2(n873), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G95), .A2(n878), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G107), .A2(n874), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n887) );
  NAND2_X1 U883 ( .A1(G1991), .A2(n887), .ZN(n801) );
  XOR2_X1 U884 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n793) );
  NAND2_X1 U885 ( .A1(G105), .A2(n878), .ZN(n792) );
  XNOR2_X1 U886 ( .A(n793), .B(n792), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G141), .A2(n877), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G129), .A2(n873), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n874), .A2(G117), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n886) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n886), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n1006) );
  NAND2_X1 U895 ( .A1(n1006), .A2(n818), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT91), .ZN(n810) );
  INV_X1 U897 ( .A(n810), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n813), .A2(n803), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n821) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n886), .ZN(n1010) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n887), .ZN(n1002) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U903 ( .A1(n1002), .A2(n808), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n1010), .A2(n811), .ZN(n812) );
  XNOR2_X1 U906 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n893), .A2(n815), .ZN(n1014) );
  NAND2_X1 U909 ( .A1(n816), .A2(n1014), .ZN(n817) );
  XOR2_X1 U910 ( .A(KEYINPUT103), .B(n817), .Z(n819) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U916 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(G188) );
  NOR2_X1 U919 ( .A1(n828), .A2(n827), .ZN(G325) );
  XNOR2_X1 U920 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  XOR2_X1 U925 ( .A(G2678), .B(KEYINPUT106), .Z(n830) );
  XNOR2_X1 U926 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT42), .B(G2090), .Z(n832) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2096), .B(G2100), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n838) );
  XOR2_X1 U934 ( .A(G2078), .B(G2084), .Z(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1961), .B(G1971), .Z(n840) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1976), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U939 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(G2474), .B(G1956), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1981), .B(G1966), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U946 ( .A(KEYINPUT113), .B(n848), .Z(n850) );
  XNOR2_X1 U947 ( .A(G171), .B(G286), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n957), .B(n942), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  NOR2_X1 U951 ( .A1(G37), .A2(n853), .ZN(G397) );
  NAND2_X1 U952 ( .A1(G100), .A2(n878), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G112), .A2(n874), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U955 ( .A(KEYINPUT108), .B(n856), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G124), .A2(n873), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U958 ( .A1(n877), .A2(G136), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U961 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G127), .A2(n873), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G115), .A2(n874), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n878), .A2(G103), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT110), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G139), .A2(n877), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n996) );
  XOR2_X1 U971 ( .A(n1001), .B(n996), .Z(n872) );
  XNOR2_X1 U972 ( .A(G160), .B(G162), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n885) );
  NAND2_X1 U974 ( .A1(G130), .A2(n873), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G118), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n883) );
  NAND2_X1 U977 ( .A1(G142), .A2(n877), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G106), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(n885), .B(n884), .Z(n895) );
  XNOR2_X1 U983 ( .A(G164), .B(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(KEYINPUT48), .Z(n891) );
  XNOR2_X1 U986 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT112), .B(n897), .ZN(G395) );
  XOR2_X1 U992 ( .A(G2443), .B(G2451), .Z(n899) );
  XNOR2_X1 U993 ( .A(G2446), .B(G2454), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n900), .B(G2427), .Z(n902) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U998 ( .A(G2435), .B(KEYINPUT104), .Z(n904) );
  XNOR2_X1 U999 ( .A(G2430), .B(G2438), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1001 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1002 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  INV_X1 U1011 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(G34), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(G2084), .B(n915), .ZN(n931) );
  XNOR2_X1 U1015 ( .A(G2090), .B(G35), .ZN(n929) );
  XOR2_X1 U1016 ( .A(G1991), .B(G25), .Z(n916) );
  NAND2_X1 U1017 ( .A1(n916), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1018 ( .A(G1996), .B(G32), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n917), .B(G27), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(KEYINPUT116), .B(n920), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G26), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(G33), .B(G2072), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n932) );
  XNOR2_X1 U1031 ( .A(n933), .B(n932), .ZN(n934) );
  INV_X1 U1032 ( .A(G29), .ZN(n1020) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n1020), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n935), .A2(G11), .ZN(n995) );
  XNOR2_X1 U1035 ( .A(G16), .B(KEYINPUT56), .ZN(n964) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n937) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT57), .ZN(n962) );
  NAND2_X1 U1039 ( .A1(G1971), .A2(G303), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(G171), .B(G1961), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(n941), .B(KEYINPUT119), .ZN(n944) );
  XOR2_X1 U1043 ( .A(G1348), .B(n942), .Z(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(KEYINPUT120), .B(n945), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n946), .B(G1956), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n947), .B(KEYINPUT121), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n956), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G1341), .B(n957), .Z(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT123), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n993) );
  INV_X1 U1058 ( .A(G16), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G5), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G1976), .B(G23), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G1986), .B(KEYINPUT127), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(n969), .B(G24), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1068 ( .A(KEYINPUT58), .B(n972), .Z(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(KEYINPUT59), .B(G1348), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(n975), .B(G4), .ZN(n984) );
  XOR2_X1 U1072 ( .A(n976), .B(G20), .Z(n982) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n977), .B(KEYINPUT124), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(G19), .B(G1341), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT125), .B(n980), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT126), .B(n985), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(KEYINPUT60), .B(n986), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT61), .B(n989), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1024) );
  XNOR2_X1 U1087 ( .A(G160), .B(G2084), .ZN(n1008) );
  XOR2_X1 U1088 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT50), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT114), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT52), .B(n1018), .Z(n1019) );
  NOR2_X1 U1104 ( .A1(KEYINPUT55), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(n1022), .B(KEYINPUT115), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

