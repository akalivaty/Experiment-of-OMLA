

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n745), .ZN(n766) );
  NOR2_X1 U553 ( .A1(G651), .A2(G543), .ZN(n687) );
  NOR2_X1 U554 ( .A1(G651), .A2(n556), .ZN(n697) );
  NAND2_X2 U555 ( .A1(n787), .A2(n786), .ZN(n795) );
  XNOR2_X2 U556 ( .A(n825), .B(KEYINPUT99), .ZN(n742) );
  NOR2_X4 U557 ( .A1(G2104), .A2(G2105), .ZN(n569) );
  NAND2_X1 U558 ( .A1(n735), .A2(n734), .ZN(n825) );
  AND2_X1 U559 ( .A1(n540), .A2(n538), .ZN(n537) );
  NOR2_X1 U560 ( .A1(n530), .A2(n526), .ZN(n525) );
  OR2_X1 U561 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U562 ( .A1(n851), .A2(G1966), .ZN(n534) );
  AND2_X1 U563 ( .A1(n613), .A2(n612), .ZN(n735) );
  NAND2_X1 U564 ( .A1(n791), .A2(n532), .ZN(n531) );
  AND2_X1 U565 ( .A1(n549), .A2(n520), .ZN(n548) );
  OR2_X1 U566 ( .A1(n968), .A2(KEYINPUT108), .ZN(n549) );
  INV_X1 U567 ( .A(KEYINPUT108), .ZN(n545) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n826) );
  NAND2_X1 U569 ( .A1(n843), .A2(n842), .ZN(n543) );
  NAND2_X1 U570 ( .A1(n570), .A2(G2104), .ZN(n571) );
  NOR2_X1 U571 ( .A1(n794), .A2(n534), .ZN(n778) );
  NOR2_X1 U572 ( .A1(n795), .A2(n531), .ZN(n530) );
  NAND2_X1 U573 ( .A1(n529), .A2(n527), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n528), .A2(KEYINPUT106), .ZN(n527) );
  OR2_X1 U575 ( .A1(G286), .A2(n531), .ZN(n529) );
  AND2_X1 U576 ( .A1(G286), .A2(KEYINPUT106), .ZN(n524) );
  NOR2_X1 U577 ( .A1(G2084), .A2(n767), .ZN(n794) );
  NAND2_X1 U578 ( .A1(n547), .A2(n544), .ZN(n552) );
  NAND2_X1 U579 ( .A1(n546), .A2(n545), .ZN(n544) );
  AND2_X1 U580 ( .A1(n550), .A2(n548), .ZN(n547) );
  NOR2_X1 U581 ( .A1(n542), .A2(n859), .ZN(n541) );
  INV_X1 U582 ( .A(n858), .ZN(n542) );
  NOR2_X1 U583 ( .A1(n858), .A2(KEYINPUT109), .ZN(n539) );
  XNOR2_X1 U584 ( .A(n616), .B(n615), .ZN(n733) );
  NOR2_X2 U585 ( .A1(G2104), .A2(n570), .ZN(n611) );
  NOR2_X1 U586 ( .A1(n851), .A2(n802), .ZN(n520) );
  AND2_X1 U587 ( .A1(n735), .A2(n553), .ZN(G160) );
  AND2_X1 U588 ( .A1(n870), .A2(n869), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n525), .A2(n523), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n795), .A2(n524), .ZN(n523) );
  INV_X1 U591 ( .A(n791), .ZN(n528) );
  INV_X1 U592 ( .A(KEYINPUT106), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n533), .A2(G8), .ZN(n793) );
  NOR2_X1 U594 ( .A1(n796), .A2(n534), .ZN(n797) );
  NAND2_X1 U595 ( .A1(n537), .A2(n535), .ZN(n871) );
  NAND2_X1 U596 ( .A1(n536), .A2(n859), .ZN(n535) );
  INV_X1 U597 ( .A(n543), .ZN(n536) );
  NOR2_X1 U598 ( .A1(n539), .A2(n522), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n543), .A2(n541), .ZN(n540) );
  INV_X1 U600 ( .A(n847), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n847), .A2(n551), .ZN(n550) );
  AND2_X1 U602 ( .A1(n968), .A2(KEYINPUT108), .ZN(n551) );
  XNOR2_X1 U603 ( .A(n552), .B(KEYINPUT64), .ZN(n804) );
  INV_X1 U604 ( .A(n733), .ZN(n553) );
  INV_X1 U605 ( .A(G2105), .ZN(n570) );
  NAND2_X1 U606 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X2 U607 ( .A(n569), .B(n568), .ZN(n929) );
  XNOR2_X1 U608 ( .A(KEYINPUT70), .B(n559), .ZN(n554) );
  AND2_X1 U609 ( .A1(G78), .A2(n688), .ZN(n555) );
  INV_X1 U610 ( .A(KEYINPUT105), .ZN(n777) );
  OR2_X2 U611 ( .A1(n776), .A2(n775), .ZN(n851) );
  INV_X1 U612 ( .A(G40), .ZN(n732) );
  NOR2_X1 U613 ( .A1(n733), .A2(n732), .ZN(n734) );
  BUF_X1 U614 ( .A(n614), .Z(n931) );
  XNOR2_X1 U615 ( .A(n623), .B(KEYINPUT13), .ZN(n624) );
  INV_X1 U616 ( .A(KEYINPUT17), .ZN(n568) );
  NAND2_X1 U617 ( .A1(n560), .A2(n554), .ZN(n561) );
  XNOR2_X1 U618 ( .A(n625), .B(n624), .ZN(n628) );
  XNOR2_X1 U619 ( .A(n571), .B(KEYINPUT65), .ZN(n614) );
  XNOR2_X1 U620 ( .A(n640), .B(n639), .ZN(n957) );
  XNOR2_X1 U621 ( .A(KEYINPUT23), .B(KEYINPUT66), .ZN(n615) );
  XOR2_X1 U622 ( .A(KEYINPUT71), .B(n564), .Z(G299) );
  XOR2_X1 U623 ( .A(G543), .B(KEYINPUT0), .Z(n556) );
  NAND2_X1 U624 ( .A1(n697), .A2(G53), .ZN(n563) );
  INV_X1 U625 ( .A(G651), .ZN(n557) );
  NOR2_X1 U626 ( .A1(n556), .A2(n557), .ZN(n688) );
  NOR2_X1 U627 ( .A1(G543), .A2(n557), .ZN(n558) );
  XOR2_X2 U628 ( .A(KEYINPUT1), .B(n558), .Z(n702) );
  NAND2_X1 U629 ( .A1(G65), .A2(n702), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n687), .A2(G91), .ZN(n559) );
  NOR2_X1 U631 ( .A1(n555), .A2(n561), .ZN(n562) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G126), .A2(n611), .ZN(n566) );
  AND2_X1 U634 ( .A1(G2104), .A2(G2105), .ZN(n925) );
  NAND2_X1 U635 ( .A1(G114), .A2(n925), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U637 ( .A(KEYINPUT92), .B(n567), .Z(n575) );
  NAND2_X1 U638 ( .A1(G138), .A2(n929), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G102), .A2(n614), .ZN(n572) );
  AND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(G164) );
  NAND2_X1 U642 ( .A1(n687), .A2(G89), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT4), .B(n576), .Z(n579) );
  NAND2_X1 U644 ( .A1(n688), .A2(G76), .ZN(n577) );
  XOR2_X1 U645 ( .A(KEYINPUT78), .B(n577), .Z(n578) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(KEYINPUT5), .B(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT79), .ZN(n587) );
  NAND2_X1 U649 ( .A1(G63), .A2(n702), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G51), .A2(n697), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n585) );
  XOR2_X1 U652 ( .A(KEYINPUT80), .B(KEYINPUT6), .Z(n584) );
  XNOR2_X1 U653 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U655 ( .A(KEYINPUT7), .B(n588), .ZN(G168) );
  XOR2_X1 U656 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U657 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U658 ( .A(G2443), .B(G2446), .Z(n590) );
  XNOR2_X1 U659 ( .A(G2427), .B(G2451), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n590), .B(n589), .ZN(n596) );
  XOR2_X1 U661 ( .A(G2430), .B(G2454), .Z(n592) );
  XNOR2_X1 U662 ( .A(G1348), .B(G1341), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n592), .B(n591), .ZN(n594) );
  XOR2_X1 U664 ( .A(G2435), .B(G2438), .Z(n593) );
  XNOR2_X1 U665 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U666 ( .A(n596), .B(n595), .Z(n597) );
  AND2_X1 U667 ( .A1(G14), .A2(n597), .ZN(G401) );
  NAND2_X1 U668 ( .A1(n688), .A2(G77), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT69), .B(n598), .Z(n600) );
  NAND2_X1 U670 ( .A1(n687), .A2(G90), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(KEYINPUT9), .B(n601), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G64), .A2(n702), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G52), .A2(n697), .ZN(n602) );
  AND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(G301) );
  INV_X1 U677 ( .A(G301), .ZN(G171) );
  AND2_X1 U678 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U679 ( .A(G132), .ZN(G219) );
  INV_X1 U680 ( .A(G82), .ZN(G220) );
  INV_X1 U681 ( .A(G57), .ZN(G237) );
  NAND2_X1 U682 ( .A1(n929), .A2(G137), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G113), .A2(n925), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  OR2_X1 U685 ( .A1(n608), .A2(KEYINPUT67), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n608), .A2(KEYINPUT67), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G125), .A2(n611), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G101), .A2(n614), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G7), .A2(G661), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U692 ( .A(G223), .ZN(n872) );
  NAND2_X1 U693 ( .A1(n872), .A2(G567), .ZN(n618) );
  XOR2_X1 U694 ( .A(KEYINPUT11), .B(n618), .Z(G234) );
  NAND2_X1 U695 ( .A1(G81), .A2(n687), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT12), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n620), .B(KEYINPUT72), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G68), .A2(n688), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n625) );
  XNOR2_X1 U700 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n702), .A2(G56), .ZN(n626) );
  XOR2_X1 U702 ( .A(KEYINPUT14), .B(n626), .Z(n627) );
  NOR2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n697), .A2(G43), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n960) );
  INV_X1 U706 ( .A(G860), .ZN(n646) );
  OR2_X1 U707 ( .A1(n960), .A2(n646), .ZN(G153) );
  INV_X1 U708 ( .A(G868), .ZN(n713) );
  NOR2_X1 U709 ( .A1(n713), .A2(G171), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(KEYINPUT75), .ZN(n642) );
  NAND2_X1 U711 ( .A1(G92), .A2(n687), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G66), .A2(n702), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U714 ( .A(KEYINPUT76), .B(n634), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G79), .A2(n688), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G54), .A2(n697), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U719 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n639) );
  OR2_X1 U720 ( .A1(G868), .A2(n957), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(G284) );
  XNOR2_X1 U722 ( .A(KEYINPUT81), .B(G868), .ZN(n643) );
  NOR2_X1 U723 ( .A1(G286), .A2(n643), .ZN(n645) );
  NOR2_X1 U724 ( .A1(G868), .A2(G299), .ZN(n644) );
  NOR2_X1 U725 ( .A1(n645), .A2(n644), .ZN(G297) );
  NAND2_X1 U726 ( .A1(n646), .A2(G559), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n647), .A2(n957), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n648), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U729 ( .A1(n957), .A2(G868), .ZN(n649) );
  XOR2_X1 U730 ( .A(KEYINPUT83), .B(n649), .Z(n650) );
  NOR2_X1 U731 ( .A1(G559), .A2(n650), .ZN(n653) );
  NOR2_X1 U732 ( .A1(G868), .A2(n960), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n651), .B(KEYINPUT82), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(G282) );
  NAND2_X1 U735 ( .A1(n611), .A2(G123), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(KEYINPUT18), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G111), .A2(n925), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G135), .A2(n929), .ZN(n658) );
  NAND2_X1 U740 ( .A1(G99), .A2(n931), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n1042) );
  XNOR2_X1 U743 ( .A(n1042), .B(G2096), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(KEYINPUT84), .ZN(n663) );
  INV_X1 U745 ( .A(G2100), .ZN(n662) );
  NAND2_X1 U746 ( .A1(n663), .A2(n662), .ZN(G156) );
  NAND2_X1 U747 ( .A1(G93), .A2(n687), .ZN(n665) );
  NAND2_X1 U748 ( .A1(G80), .A2(n688), .ZN(n664) );
  NAND2_X1 U749 ( .A1(n665), .A2(n664), .ZN(n669) );
  NAND2_X1 U750 ( .A1(G67), .A2(n702), .ZN(n667) );
  NAND2_X1 U751 ( .A1(G55), .A2(n697), .ZN(n666) );
  NAND2_X1 U752 ( .A1(n667), .A2(n666), .ZN(n668) );
  OR2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n714) );
  NAND2_X1 U754 ( .A1(G559), .A2(n957), .ZN(n670) );
  XOR2_X1 U755 ( .A(n960), .B(n670), .Z(n710) );
  XNOR2_X1 U756 ( .A(KEYINPUT85), .B(n710), .ZN(n671) );
  NOR2_X1 U757 ( .A1(G860), .A2(n671), .ZN(n672) );
  XOR2_X1 U758 ( .A(n714), .B(n672), .Z(G145) );
  NAND2_X1 U759 ( .A1(G86), .A2(n687), .ZN(n674) );
  NAND2_X1 U760 ( .A1(G61), .A2(n702), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n688), .A2(G73), .ZN(n675) );
  XOR2_X1 U763 ( .A(KEYINPUT2), .B(n675), .Z(n676) );
  NOR2_X1 U764 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n697), .A2(G48), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(G305) );
  NAND2_X1 U767 ( .A1(G85), .A2(n687), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G72), .A2(n688), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G60), .A2(n702), .ZN(n683) );
  NAND2_X1 U771 ( .A1(G47), .A2(n697), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U774 ( .A(KEYINPUT68), .B(n686), .Z(G290) );
  NAND2_X1 U775 ( .A1(G62), .A2(n702), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G88), .A2(n687), .ZN(n690) );
  NAND2_X1 U777 ( .A1(G75), .A2(n688), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U779 ( .A1(G50), .A2(n697), .ZN(n691) );
  XNOR2_X1 U780 ( .A(KEYINPUT87), .B(n691), .ZN(n692) );
  NOR2_X1 U781 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U783 ( .A(n696), .B(KEYINPUT88), .ZN(G303) );
  NAND2_X1 U784 ( .A1(G49), .A2(n697), .ZN(n699) );
  NAND2_X1 U785 ( .A1(G74), .A2(G651), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U787 ( .A(KEYINPUT86), .B(n700), .ZN(n701) );
  NOR2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n556), .A2(G87), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n704), .A2(n703), .ZN(G288) );
  XOR2_X1 U791 ( .A(G290), .B(n714), .Z(n705) );
  XNOR2_X1 U792 ( .A(n705), .B(KEYINPUT19), .ZN(n706) );
  XNOR2_X1 U793 ( .A(G305), .B(n706), .ZN(n708) );
  INV_X1 U794 ( .A(G299), .ZN(n964) );
  XNOR2_X1 U795 ( .A(n964), .B(G303), .ZN(n707) );
  XNOR2_X1 U796 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U797 ( .A(n709), .B(G288), .ZN(n940) );
  XNOR2_X1 U798 ( .A(n940), .B(n710), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n711), .A2(G868), .ZN(n712) );
  XOR2_X1 U800 ( .A(KEYINPUT89), .B(n712), .Z(n716) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n716), .A2(n715), .ZN(G295) );
  XOR2_X1 U803 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n718) );
  NAND2_X1 U804 ( .A1(G2078), .A2(G2084), .ZN(n717) );
  XNOR2_X1 U805 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U806 ( .A1(G2090), .A2(n719), .ZN(n720) );
  XNOR2_X1 U807 ( .A(KEYINPUT21), .B(n720), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n721), .A2(G2072), .ZN(G158) );
  NAND2_X1 U809 ( .A1(G69), .A2(G120), .ZN(n722) );
  NOR2_X1 U810 ( .A1(G237), .A2(n722), .ZN(n723) );
  NAND2_X1 U811 ( .A1(G108), .A2(n723), .ZN(n876) );
  NAND2_X1 U812 ( .A1(G567), .A2(n876), .ZN(n724) );
  XNOR2_X1 U813 ( .A(n724), .B(KEYINPUT91), .ZN(n729) );
  NOR2_X1 U814 ( .A1(G220), .A2(G219), .ZN(n725) );
  XNOR2_X1 U815 ( .A(KEYINPUT22), .B(n725), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n726), .A2(G96), .ZN(n727) );
  OR2_X1 U817 ( .A1(G218), .A2(n727), .ZN(n877) );
  AND2_X1 U818 ( .A1(G2106), .A2(n877), .ZN(n728) );
  NOR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(G319) );
  INV_X1 U820 ( .A(G319), .ZN(n731) );
  NAND2_X1 U821 ( .A1(G483), .A2(G661), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n875) );
  NAND2_X1 U823 ( .A1(n875), .A2(G36), .ZN(G176) );
  AND2_X1 U824 ( .A1(n826), .A2(G2072), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n742), .A2(n736), .ZN(n737) );
  XNOR2_X1 U826 ( .A(n737), .B(KEYINPUT27), .ZN(n739) );
  INV_X1 U827 ( .A(G1956), .ZN(n1001) );
  NAND2_X1 U828 ( .A1(n742), .A2(n826), .ZN(n745) );
  INV_X1 U829 ( .A(n745), .ZN(n775) );
  NOR2_X1 U830 ( .A1(n1001), .A2(n775), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n760) );
  NOR2_X1 U832 ( .A1(n964), .A2(n760), .ZN(n740) );
  XOR2_X1 U833 ( .A(n740), .B(KEYINPUT28), .Z(n759) );
  AND2_X1 U834 ( .A1(n826), .A2(G1996), .ZN(n741) );
  AND2_X1 U835 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n743), .B(KEYINPUT26), .ZN(n744) );
  INV_X1 U837 ( .A(n744), .ZN(n747) );
  INV_X1 U838 ( .A(n766), .ZN(n767) );
  NAND2_X1 U839 ( .A1(n767), .A2(G1341), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n960), .A2(n748), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n957), .A2(n751), .ZN(n749) );
  XNOR2_X1 U843 ( .A(n749), .B(KEYINPUT103), .ZN(n750) );
  AND2_X1 U844 ( .A1(n759), .A2(n750), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n957), .A2(n751), .ZN(n752) );
  XNOR2_X1 U846 ( .A(n752), .B(KEYINPUT102), .ZN(n756) );
  NOR2_X1 U847 ( .A1(n775), .A2(G1348), .ZN(n754) );
  NOR2_X1 U848 ( .A1(G2067), .A2(n767), .ZN(n753) );
  NOR2_X1 U849 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n764) );
  INV_X1 U852 ( .A(n759), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n964), .A2(n760), .ZN(n761) );
  XNOR2_X1 U854 ( .A(n765), .B(KEYINPUT29), .ZN(n773) );
  OR2_X1 U855 ( .A1(n766), .A2(G1961), .ZN(n770) );
  XNOR2_X1 U856 ( .A(G2078), .B(KEYINPUT25), .ZN(n768) );
  XNOR2_X1 U857 ( .A(n768), .B(KEYINPUT100), .ZN(n984) );
  NAND2_X1 U858 ( .A1(n766), .A2(n984), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n782) );
  AND2_X1 U860 ( .A1(n782), .A2(G171), .ZN(n771) );
  XNOR2_X1 U861 ( .A(KEYINPUT101), .B(n771), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT104), .ZN(n787) );
  INV_X1 U864 ( .A(G8), .ZN(n776) );
  XNOR2_X1 U865 ( .A(n778), .B(n777), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n779), .A2(G8), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT30), .B(n780), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n781), .A2(G168), .ZN(n784) );
  NOR2_X1 U869 ( .A1(G171), .A2(n782), .ZN(n783) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U871 ( .A(KEYINPUT31), .B(n785), .Z(n786) );
  NOR2_X1 U872 ( .A1(G1971), .A2(n851), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G2090), .A2(n767), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n790), .A2(G303), .ZN(n791) );
  XOR2_X1 U876 ( .A(KEYINPUT107), .B(KEYINPUT32), .Z(n792) );
  XNOR2_X1 U877 ( .A(n793), .B(n792), .ZN(n800) );
  NAND2_X1 U878 ( .A1(G8), .A2(n794), .ZN(n798) );
  INV_X1 U879 ( .A(n795), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U881 ( .A1(n800), .A2(n799), .ZN(n847) );
  NOR2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n805) );
  NOR2_X1 U883 ( .A1(G303), .A2(G1971), .ZN(n801) );
  NOR2_X1 U884 ( .A1(n805), .A2(n801), .ZN(n968) );
  NAND2_X1 U885 ( .A1(G1976), .A2(G288), .ZN(n967) );
  INV_X1 U886 ( .A(n967), .ZN(n802) );
  INV_X1 U887 ( .A(KEYINPUT33), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n843) );
  NAND2_X1 U889 ( .A1(n805), .A2(KEYINPUT33), .ZN(n806) );
  NOR2_X1 U890 ( .A1(n806), .A2(n851), .ZN(n841) );
  XOR2_X1 U891 ( .A(G1981), .B(G305), .Z(n953) );
  NAND2_X1 U892 ( .A1(n925), .A2(G107), .ZN(n807) );
  XOR2_X1 U893 ( .A(KEYINPUT93), .B(n807), .Z(n809) );
  NAND2_X1 U894 ( .A1(n611), .A2(G119), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U896 ( .A(KEYINPUT94), .B(n810), .Z(n814) );
  NAND2_X1 U897 ( .A1(G131), .A2(n929), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G95), .A2(n931), .ZN(n811) );
  AND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n921) );
  AND2_X1 U901 ( .A1(n921), .A2(G1991), .ZN(n824) );
  NAND2_X1 U902 ( .A1(G105), .A2(n931), .ZN(n815) );
  XOR2_X1 U903 ( .A(KEYINPUT38), .B(n815), .Z(n820) );
  NAND2_X1 U904 ( .A1(G129), .A2(n611), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G117), .A2(n925), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U907 ( .A(KEYINPUT95), .B(n818), .Z(n819) );
  NOR2_X1 U908 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n929), .A2(G141), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(n910) );
  AND2_X1 U911 ( .A1(n910), .A2(G1996), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n1038) );
  NOR2_X1 U913 ( .A1(n826), .A2(n825), .ZN(n869) );
  XOR2_X1 U914 ( .A(n869), .B(KEYINPUT96), .Z(n827) );
  NOR2_X1 U915 ( .A1(n1038), .A2(n827), .ZN(n862) );
  XNOR2_X1 U916 ( .A(KEYINPUT97), .B(n862), .ZN(n837) );
  XNOR2_X1 U917 ( .A(G2067), .B(KEYINPUT37), .ZN(n867) );
  NAND2_X1 U918 ( .A1(G140), .A2(n929), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G104), .A2(n931), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U921 ( .A(KEYINPUT34), .B(n830), .ZN(n835) );
  NAND2_X1 U922 ( .A1(G128), .A2(n611), .ZN(n832) );
  NAND2_X1 U923 ( .A1(G116), .A2(n925), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U925 ( .A(KEYINPUT35), .B(n833), .Z(n834) );
  NOR2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U927 ( .A(KEYINPUT36), .B(n836), .ZN(n906) );
  NOR2_X1 U928 ( .A1(n867), .A2(n906), .ZN(n1041) );
  NAND2_X1 U929 ( .A1(n869), .A2(n1041), .ZN(n865) );
  NAND2_X1 U930 ( .A1(n837), .A2(n865), .ZN(n838) );
  XOR2_X1 U931 ( .A(n838), .B(KEYINPUT98), .Z(n855) );
  AND2_X1 U932 ( .A1(n953), .A2(n855), .ZN(n839) );
  XNOR2_X1 U933 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U934 ( .A1(n869), .A2(n959), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n839), .A2(n844), .ZN(n840) );
  NOR2_X1 U936 ( .A1(n841), .A2(n840), .ZN(n842) );
  INV_X1 U937 ( .A(n844), .ZN(n857) );
  NOR2_X1 U938 ( .A1(G2090), .A2(G303), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G8), .A2(n845), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n851), .A2(n848), .ZN(n853) );
  NOR2_X1 U942 ( .A1(G1981), .A2(G305), .ZN(n849) );
  XOR2_X1 U943 ( .A(n849), .B(KEYINPUT24), .Z(n850) );
  OR2_X1 U944 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U945 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U946 ( .A1(n855), .A2(n854), .ZN(n856) );
  OR2_X1 U947 ( .A1(n857), .A2(n856), .ZN(n858) );
  INV_X1 U948 ( .A(KEYINPUT109), .ZN(n859) );
  NOR2_X1 U949 ( .A1(G1996), .A2(n910), .ZN(n1034) );
  NOR2_X1 U950 ( .A1(G1991), .A2(n921), .ZN(n1043) );
  NOR2_X1 U951 ( .A1(G1986), .A2(G290), .ZN(n860) );
  NOR2_X1 U952 ( .A1(n1043), .A2(n860), .ZN(n861) );
  NOR2_X1 U953 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U954 ( .A1(n1034), .A2(n863), .ZN(n864) );
  XNOR2_X1 U955 ( .A(KEYINPUT39), .B(n864), .ZN(n866) );
  NAND2_X1 U956 ( .A1(n866), .A2(n865), .ZN(n868) );
  NAND2_X1 U957 ( .A1(n867), .A2(n906), .ZN(n1047) );
  NAND2_X1 U958 ( .A1(n868), .A2(n1047), .ZN(n870) );
  XNOR2_X1 U959 ( .A(n871), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U960 ( .A1(G2106), .A2(n872), .ZN(G217) );
  AND2_X1 U961 ( .A1(G15), .A2(G2), .ZN(n873) );
  NAND2_X1 U962 ( .A1(G661), .A2(n873), .ZN(G259) );
  NAND2_X1 U963 ( .A1(G3), .A2(G1), .ZN(n874) );
  NAND2_X1 U964 ( .A1(n875), .A2(n874), .ZN(G188) );
  INV_X1 U966 ( .A(G120), .ZN(G236) );
  INV_X1 U967 ( .A(G96), .ZN(G221) );
  INV_X1 U968 ( .A(G69), .ZN(G235) );
  NOR2_X1 U969 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U970 ( .A(KEYINPUT110), .B(n878), .ZN(G325) );
  INV_X1 U971 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U972 ( .A(G1976), .B(KEYINPUT41), .ZN(n888) );
  XOR2_X1 U973 ( .A(G1971), .B(G1956), .Z(n880) );
  XNOR2_X1 U974 ( .A(G1986), .B(G1966), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U976 ( .A(G1981), .B(G1961), .Z(n882) );
  XNOR2_X1 U977 ( .A(G1996), .B(G1991), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U979 ( .A(n884), .B(n883), .Z(n886) );
  XNOR2_X1 U980 ( .A(KEYINPUT112), .B(G2474), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n888), .B(n887), .ZN(G229) );
  XOR2_X1 U983 ( .A(KEYINPUT111), .B(G2090), .Z(n890) );
  XNOR2_X1 U984 ( .A(G2078), .B(G2072), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U986 ( .A(n891), .B(G2100), .Z(n893) );
  XNOR2_X1 U987 ( .A(G2067), .B(G2084), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U989 ( .A(G2096), .B(G2678), .Z(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U992 ( .A(n897), .B(n896), .Z(G227) );
  NAND2_X1 U993 ( .A1(G112), .A2(n925), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G100), .A2(n931), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n900), .B(KEYINPUT113), .ZN(n902) );
  NAND2_X1 U997 ( .A1(G136), .A2(n929), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n611), .A2(G124), .ZN(n903) );
  XOR2_X1 U1000 ( .A(KEYINPUT44), .B(n903), .Z(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(G162) );
  XNOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n906), .B(n1042), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(n909), .B(G162), .Z(n912) );
  XOR2_X1 U1006 ( .A(G160), .B(n910), .Z(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n920) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n929), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(G103), .A2(n931), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(G127), .A2(n611), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(G115), .A2(n925), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1014 ( .A(KEYINPUT47), .B(n917), .Z(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n1029) );
  XOR2_X1 U1016 ( .A(n920), .B(n1029), .Z(n923) );
  XOR2_X1 U1017 ( .A(G164), .B(n921), .Z(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n938) );
  NAND2_X1 U1019 ( .A1(n611), .A2(G130), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(KEYINPUT114), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(G118), .A2(n925), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1023 ( .A(KEYINPUT115), .B(n928), .Z(n936) );
  NAND2_X1 U1024 ( .A1(n929), .A2(G142), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(n930), .B(KEYINPUT116), .ZN(n933) );
  NAND2_X1 U1026 ( .A1(G106), .A2(n931), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1028 ( .A(KEYINPUT45), .B(n934), .Z(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(n938), .B(n937), .ZN(n939) );
  NOR2_X1 U1031 ( .A1(G37), .A2(n939), .ZN(G395) );
  XNOR2_X1 U1032 ( .A(n960), .B(n940), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G171), .B(n957), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n942), .B(n941), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G286), .B(n943), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(G37), .A2(n944), .ZN(G397) );
  XNOR2_X1 U1037 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(G229), .A2(G227), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n946), .B(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(G319), .A2(n947), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(G401), .A2(n948), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT118), .B(n949), .ZN(n951) );
  NOR2_X1 U1043 ( .A1(G395), .A2(G397), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(G225) );
  INV_X1 U1045 ( .A(G225), .ZN(G308) );
  INV_X1 U1046 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1047 ( .A(G16), .B(KEYINPUT56), .Z(n980) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n952), .B(KEYINPUT120), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n955) );
  XNOR2_X1 U1052 ( .A(n956), .B(n955), .ZN(n975) );
  XOR2_X1 U1053 ( .A(G1348), .B(n957), .Z(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G1341), .B(KEYINPUT123), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n973) );
  XNOR2_X1 U1058 ( .A(n964), .B(G1956), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(G1971), .A2(G303), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1063 ( .A(KEYINPUT122), .B(n971), .Z(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G1961), .B(G301), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(KEYINPUT124), .B(n978), .ZN(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n1058) );
  XNOR2_X1 U1070 ( .A(G2090), .B(G35), .ZN(n993) );
  XOR2_X1 U1071 ( .A(G2067), .B(G26), .Z(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(G28), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G1991), .B(G25), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G2072), .B(G33), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n988) );
  XOR2_X1 U1076 ( .A(n984), .B(G27), .Z(n986) );
  XNOR2_X1 U1077 ( .A(G1996), .B(G32), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n991), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1083 ( .A(G2084), .B(G34), .Z(n994) );
  XNOR2_X1 U1084 ( .A(KEYINPUT54), .B(n994), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(G29), .A2(KEYINPUT55), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n997), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(G11), .A2(n998), .ZN(n1028) );
  INV_X1 U1089 ( .A(KEYINPUT55), .ZN(n1052) );
  OR2_X1 U1090 ( .A1(n1052), .A2(n999), .ZN(n1026) );
  XNOR2_X1 U1091 ( .A(G5), .B(G1961), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT125), .ZN(n1013) );
  XNOR2_X1 U1093 ( .A(G20), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1006) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1019) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1017) );
  XNOR2_X1 U1107 ( .A(G1971), .B(G22), .ZN(n1015) );
  XNOR2_X1 U1108 ( .A(G23), .B(G1976), .ZN(n1014) );
  NOR2_X1 U1109 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1110 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1111 ( .A(n1019), .B(n1018), .Z(n1020) );
  NOR2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1022), .ZN(n1024) );
  INV_X1 U1114 ( .A(G16), .ZN(n1023) );
  NAND2_X1 U1115 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1056) );
  XOR2_X1 U1118 ( .A(G2072), .B(n1029), .Z(n1031) );
  XOR2_X1 U1119 ( .A(G164), .B(G2078), .Z(n1030) );
  NOR2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1121 ( .A(KEYINPUT50), .B(n1032), .ZN(n1037) );
  XOR2_X1 U1122 ( .A(G2090), .B(G162), .Z(n1033) );
  NOR2_X1 U1123 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1124 ( .A(KEYINPUT51), .B(n1035), .Z(n1036) );
  NAND2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1050) );
  XNOR2_X1 U1126 ( .A(G160), .B(G2084), .ZN(n1039) );
  NAND2_X1 U1127 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1128 ( .A1(n1041), .A2(n1040), .ZN(n1045) );
  NOR2_X1 U1129 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1130 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XNOR2_X1 U1131 ( .A(KEYINPUT119), .B(n1046), .ZN(n1048) );
  NAND2_X1 U1132 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NOR2_X1 U1133 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XNOR2_X1 U1134 ( .A(KEYINPUT52), .B(n1051), .ZN(n1053) );
  NAND2_X1 U1135 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  NAND2_X1 U1136 ( .A1(n1054), .A2(G29), .ZN(n1055) );
  NAND2_X1 U1137 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  NOR2_X1 U1138 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XOR2_X1 U1139 ( .A(KEYINPUT127), .B(n1059), .Z(n1060) );
  XNOR2_X1 U1140 ( .A(KEYINPUT62), .B(n1060), .ZN(G311) );
  INV_X1 U1141 ( .A(G311), .ZN(G150) );
  INV_X1 U1142 ( .A(G303), .ZN(G166) );
endmodule

