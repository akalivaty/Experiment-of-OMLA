

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U558 ( .A1(n751), .A2(n749), .ZN(n728) );
  AND2_X1 U559 ( .A1(n745), .A2(n744), .ZN(n748) );
  INV_X1 U560 ( .A(n523), .ZN(n524) );
  NOR2_X4 U561 ( .A1(n530), .A2(n529), .ZN(n888) );
  INV_X1 U562 ( .A(n883), .ZN(n523) );
  XOR2_X2 U563 ( .A(KEYINPUT17), .B(n528), .Z(n882) );
  NOR2_X1 U564 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U565 ( .A1(n1001), .A2(n693), .ZN(n694) );
  NOR2_X1 U566 ( .A1(n717), .A2(n961), .ZN(n689) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n766) );
  NOR2_X1 U568 ( .A1(n703), .A2(n702), .ZN(n709) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U570 ( .A(n536), .B(n535), .ZN(n539) );
  NOR2_X1 U571 ( .A1(n826), .A2(n760), .ZN(n525) );
  XNOR2_X1 U572 ( .A(n746), .B(KEYINPUT104), .ZN(n747) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(KEYINPUT23), .ZN(n535) );
  AND2_X1 U574 ( .A1(n530), .A2(n529), .ZN(n883) );
  NOR2_X1 U575 ( .A1(G651), .A2(n634), .ZN(n653) );
  NOR2_X1 U576 ( .A1(n544), .A2(n543), .ZN(n687) );
  BUF_X1 U577 ( .A(n687), .Z(G160) );
  XNOR2_X2 U578 ( .A(G2104), .B(KEYINPUT66), .ZN(n530) );
  INV_X1 U579 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U580 ( .A1(G102), .A2(n524), .ZN(n527) );
  AND2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U582 ( .A1(G114), .A2(n886), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G138), .A2(n882), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G126), .A2(n888), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U588 ( .A1(G101), .A2(n883), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n888), .A2(G125), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n537), .B(KEYINPUT67), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U592 ( .A(n540), .B(KEYINPUT69), .ZN(n544) );
  NAND2_X1 U593 ( .A1(G137), .A2(n882), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G113), .A2(n886), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G57), .ZN(G237) );
  INV_X1 U598 ( .A(G132), .ZN(G219) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  XOR2_X1 U600 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  NAND2_X1 U601 ( .A1(G52), .A2(n653), .ZN(n548) );
  INV_X1 U602 ( .A(G651), .ZN(n549) );
  NOR2_X1 U603 ( .A1(G543), .A2(n549), .ZN(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT1), .B(KEYINPUT71), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n546), .B(n545), .ZN(n656) );
  NAND2_X1 U606 ( .A1(G64), .A2(n656), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n555) );
  NOR2_X1 U608 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U609 ( .A1(G90), .A2(n652), .ZN(n552) );
  OR2_X1 U610 ( .A1(n549), .A2(n634), .ZN(n550) );
  XOR2_X1 U611 ( .A(KEYINPUT70), .B(n550), .Z(n660) );
  NAND2_X1 U612 ( .A1(G77), .A2(n660), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U615 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U616 ( .A1(n652), .A2(G89), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G76), .A2(n660), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n559), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U621 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n653), .A2(G51), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n560), .B(KEYINPUT78), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G63), .A2(n656), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U632 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n570) );
  INV_X1 U633 ( .A(G223), .ZN(n839) );
  NAND2_X1 U634 ( .A1(G567), .A2(n839), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G234) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(KEYINPUT75), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n652), .A2(G81), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G68), .A2(n660), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n656), .A2(G56), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n576), .Z(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n653), .A2(G43), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n1001) );
  INV_X1 U647 ( .A(G860), .ZN(n601) );
  OR2_X1 U648 ( .A1(n1001), .A2(n601), .ZN(G153) );
  NAND2_X1 U649 ( .A1(G868), .A2(G171), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G54), .A2(n653), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G79), .A2(n660), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U653 ( .A(KEYINPUT76), .B(n583), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G92), .A2(n652), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G66), .A2(n656), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n588), .Z(n695) );
  BUF_X1 U659 ( .A(n695), .Z(n988) );
  INV_X1 U660 ( .A(G868), .ZN(n672) );
  NAND2_X1 U661 ( .A1(n988), .A2(n672), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT77), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G53), .A2(n653), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G65), .A2(n656), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U667 ( .A(KEYINPUT73), .B(n594), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n660), .A2(G78), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G91), .A2(n652), .ZN(n595) );
  AND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U673 ( .A1(G286), .A2(n672), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n602), .A2(n988), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U678 ( .A1(n988), .A2(G868), .ZN(n604) );
  XNOR2_X1 U679 ( .A(KEYINPUT80), .B(n604), .ZN(n605) );
  NOR2_X1 U680 ( .A1(G559), .A2(n605), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT81), .B(n606), .Z(n608) );
  NOR2_X1 U682 ( .A1(G868), .A2(n1001), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT82), .B(n609), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G135), .A2(n882), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G111), .A2(n886), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G123), .A2(n888), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n524), .A2(G99), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n938) );
  XNOR2_X1 U693 ( .A(n938), .B(G2096), .ZN(n618) );
  INV_X1 U694 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G559), .A2(n988), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT83), .ZN(n669) );
  XOR2_X1 U698 ( .A(n1001), .B(n669), .Z(n620) );
  NOR2_X1 U699 ( .A1(G860), .A2(n620), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G55), .A2(n653), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G67), .A2(n656), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT84), .B(n623), .Z(n627) );
  NAND2_X1 U704 ( .A1(n660), .A2(G80), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G93), .A2(n652), .ZN(n624) );
  AND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n671) );
  XNOR2_X1 U708 ( .A(n628), .B(n671), .ZN(n629) );
  XNOR2_X1 U709 ( .A(KEYINPUT85), .B(n629), .ZN(G145) );
  NAND2_X1 U710 ( .A1(G49), .A2(n653), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U713 ( .A(KEYINPUT86), .B(n632), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n656), .A2(n633), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G88), .A2(n652), .ZN(n638) );
  NAND2_X1 U718 ( .A1(G62), .A2(n656), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n660), .A2(G75), .ZN(n639) );
  XOR2_X1 U721 ( .A(KEYINPUT88), .B(n639), .Z(n640) );
  NOR2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n653), .A2(G50), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U725 ( .A(G303), .ZN(G166) );
  NAND2_X1 U726 ( .A1(G86), .A2(n652), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G61), .A2(n656), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G73), .A2(n660), .ZN(n646) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U732 ( .A(KEYINPUT87), .B(n649), .Z(n651) );
  NAND2_X1 U733 ( .A1(n653), .A2(G48), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G85), .A2(n652), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G47), .A2(n653), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n656), .A2(G60), .ZN(n657) );
  XOR2_X1 U739 ( .A(KEYINPUT72), .B(n657), .Z(n658) );
  NOR2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G72), .A2(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(G290) );
  XOR2_X1 U743 ( .A(G288), .B(n671), .Z(n664) );
  INV_X1 U744 ( .A(G299), .ZN(n710) );
  XNOR2_X1 U745 ( .A(n710), .B(G166), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G305), .ZN(n668) );
  XOR2_X1 U748 ( .A(KEYINPUT19), .B(G290), .Z(n666) );
  XNOR2_X1 U749 ( .A(n1001), .B(n666), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n668), .B(n667), .ZN(n905) );
  XNOR2_X1 U751 ( .A(n669), .B(n905), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U763 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G96), .A2(n681), .ZN(n843) );
  NAND2_X1 U765 ( .A1(n843), .A2(G2106), .ZN(n685) );
  NAND2_X1 U766 ( .A1(G69), .A2(G120), .ZN(n682) );
  NOR2_X1 U767 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U768 ( .A1(G108), .A2(n683), .ZN(n844) );
  NAND2_X1 U769 ( .A1(n844), .A2(G567), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n845) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U772 ( .A1(n845), .A2(n686), .ZN(n842) );
  NAND2_X1 U773 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G171), .ZN(G301) );
  INV_X1 U775 ( .A(n766), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n687), .A2(G40), .ZN(n767) );
  OR2_X2 U777 ( .A1(n690), .A2(n767), .ZN(n717) );
  INV_X1 U778 ( .A(G1996), .ZN(n961) );
  XOR2_X1 U779 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n688) );
  XNOR2_X1 U780 ( .A(n689), .B(n688), .ZN(n692) );
  NOR2_X1 U781 ( .A1(n690), .A2(n767), .ZN(n720) );
  NAND2_X1 U782 ( .A1(n717), .A2(G1341), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n694), .B(KEYINPUT65), .ZN(n699) );
  INV_X1 U785 ( .A(n695), .ZN(n700) );
  XNOR2_X1 U786 ( .A(n717), .B(KEYINPUT99), .ZN(n705) );
  NAND2_X1 U787 ( .A1(G2067), .A2(n705), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n717), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n701) );
  AND2_X1 U790 ( .A1(n700), .A2(n701), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n705), .A2(G2072), .ZN(n704) );
  XNOR2_X1 U794 ( .A(n704), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U795 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U796 ( .A1(n1008), .A2(n705), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n711), .A2(n710), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n715) );
  INV_X1 U799 ( .A(KEYINPUT28), .ZN(n712) );
  XNOR2_X1 U800 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U802 ( .A(n716), .B(KEYINPUT29), .ZN(n724) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n959) );
  XOR2_X1 U804 ( .A(n717), .B(KEYINPUT99), .Z(n718) );
  NOR2_X1 U805 ( .A1(n959), .A2(n718), .ZN(n719) );
  XNOR2_X1 U806 ( .A(n719), .B(KEYINPUT100), .ZN(n722) );
  NOR2_X1 U807 ( .A1(n720), .A2(G1961), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U809 ( .A1(G301), .A2(n725), .ZN(n723) );
  NOR2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n735) );
  NAND2_X1 U811 ( .A1(n725), .A2(G301), .ZN(n726) );
  XNOR2_X1 U812 ( .A(n726), .B(KEYINPUT101), .ZN(n732) );
  NAND2_X1 U813 ( .A1(G8), .A2(n717), .ZN(n826) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n826), .ZN(n751) );
  NOR2_X1 U815 ( .A1(n717), .A2(G2084), .ZN(n727) );
  XNOR2_X1 U816 ( .A(n727), .B(KEYINPUT98), .ZN(n749) );
  NAND2_X1 U817 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n730), .A2(G168), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n733), .B(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U823 ( .A(n736), .B(KEYINPUT102), .ZN(n750) );
  INV_X1 U824 ( .A(n750), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n737), .A2(G286), .ZN(n745) );
  INV_X1 U826 ( .A(G8), .ZN(n743) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n826), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n717), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U830 ( .A(KEYINPUT103), .B(n740), .Z(n741) );
  NAND2_X1 U831 ( .A1(n741), .A2(G303), .ZN(n742) );
  OR2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U833 ( .A(KEYINPUT32), .B(KEYINPUT105), .Z(n746) );
  XNOR2_X1 U834 ( .A(n748), .B(n747), .ZN(n755) );
  NAND2_X1 U835 ( .A1(n749), .A2(G8), .ZN(n753) );
  NOR2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n755), .A2(n754), .ZN(n822) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n992), .A2(n756), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n822), .A2(n757), .ZN(n758) );
  XNOR2_X1 U843 ( .A(n758), .B(KEYINPUT106), .ZN(n761) );
  NAND2_X1 U844 ( .A1(G288), .A2(G1976), .ZN(n759) );
  XOR2_X1 U845 ( .A(KEYINPUT107), .B(n759), .Z(n993) );
  INV_X1 U846 ( .A(n993), .ZN(n760) );
  AND2_X1 U847 ( .A1(n761), .A2(n525), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n762), .A2(KEYINPUT33), .ZN(n764) );
  INV_X1 U849 ( .A(KEYINPUT108), .ZN(n763) );
  XNOR2_X1 U850 ( .A(n764), .B(n763), .ZN(n819) );
  NAND2_X1 U851 ( .A1(n992), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n826), .A2(n765), .ZN(n817) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n980) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n810) );
  XNOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .ZN(n768) );
  XNOR2_X1 U856 ( .A(n768), .B(KEYINPUT90), .ZN(n781) );
  NAND2_X1 U857 ( .A1(n524), .A2(G104), .ZN(n769) );
  XOR2_X1 U858 ( .A(KEYINPUT91), .B(n769), .Z(n771) );
  NAND2_X1 U859 ( .A1(n882), .A2(G140), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n772), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G116), .A2(n886), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G128), .A2(n888), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  XNOR2_X1 U866 ( .A(KEYINPUT92), .B(n776), .ZN(n777) );
  NOR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U868 ( .A(n779), .B(KEYINPUT36), .Z(n780) );
  XNOR2_X1 U869 ( .A(KEYINPUT93), .B(n780), .ZN(n902) );
  NOR2_X1 U870 ( .A1(n781), .A2(n902), .ZN(n936) );
  NAND2_X1 U871 ( .A1(n810), .A2(n936), .ZN(n831) );
  AND2_X1 U872 ( .A1(n980), .A2(n831), .ZN(n815) );
  NAND2_X1 U873 ( .A1(n781), .A2(n902), .ZN(n935) );
  NAND2_X1 U874 ( .A1(G141), .A2(n882), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G117), .A2(n886), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n524), .A2(G105), .ZN(n784) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n888), .A2(G129), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n897) );
  NOR2_X1 U882 ( .A1(G1996), .A2(n897), .ZN(n929) );
  NAND2_X1 U883 ( .A1(G95), .A2(n524), .ZN(n789) );
  XOR2_X1 U884 ( .A(KEYINPUT96), .B(n789), .Z(n795) );
  NAND2_X1 U885 ( .A1(n888), .A2(G119), .ZN(n790) );
  XNOR2_X1 U886 ( .A(n790), .B(KEYINPUT94), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G107), .A2(n886), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U889 ( .A(KEYINPUT95), .B(n793), .Z(n794) );
  NOR2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n882), .A2(G131), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n871) );
  AND2_X1 U893 ( .A1(n871), .A2(G1991), .ZN(n799) );
  AND2_X1 U894 ( .A1(G1996), .A2(n897), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n941) );
  INV_X1 U896 ( .A(n810), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n941), .A2(n800), .ZN(n809) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n871), .ZN(n939) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U900 ( .A1(n939), .A2(n801), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n809), .A2(n802), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n929), .A2(n803), .ZN(n804) );
  XNOR2_X1 U903 ( .A(n804), .B(KEYINPUT39), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n805), .A2(n831), .ZN(n806) );
  XOR2_X1 U905 ( .A(KEYINPUT109), .B(n806), .Z(n807) );
  NAND2_X1 U906 ( .A1(n935), .A2(n807), .ZN(n808) );
  AND2_X1 U907 ( .A1(n808), .A2(n810), .ZN(n832) );
  INV_X1 U908 ( .A(n809), .ZN(n813) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U910 ( .A1(n984), .A2(n810), .ZN(n811) );
  XOR2_X1 U911 ( .A(KEYINPUT89), .B(n811), .Z(n812) );
  AND2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U913 ( .A1(n832), .A2(n814), .ZN(n835) );
  NAND2_X1 U914 ( .A1(n815), .A2(n835), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n837) );
  NOR2_X1 U917 ( .A1(G2090), .A2(G303), .ZN(n820) );
  NAND2_X1 U918 ( .A1(G8), .A2(n820), .ZN(n821) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n823), .A2(n826), .ZN(n829) );
  NOR2_X1 U921 ( .A1(G1981), .A2(G305), .ZN(n824) );
  XNOR2_X1 U922 ( .A(n824), .B(KEYINPUT24), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n825), .B(KEYINPUT97), .ZN(n827) );
  OR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  AND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n833) );
  OR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U930 ( .A(n838), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U933 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  INV_X1 U942 ( .A(n845), .ZN(G319) );
  XOR2_X1 U943 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U952 ( .A(G1971), .B(G1966), .Z(n855) );
  XNOR2_X1 U953 ( .A(G1961), .B(G1956), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(G1976), .B(G1986), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(G2474), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U961 ( .A(G1981), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G136), .A2(n882), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G112), .A2(n886), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G124), .A2(n888), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n524), .A2(G100), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(G162) );
  XOR2_X1 U971 ( .A(G160), .B(n871), .Z(n901) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n873) );
  XNOR2_X1 U973 ( .A(G164), .B(n938), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n896) );
  NAND2_X1 U975 ( .A1(G142), .A2(n882), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G106), .A2(n524), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT45), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G118), .A2(n886), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G130), .A2(n888), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n879), .Z(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n894) );
  NAND2_X1 U984 ( .A1(G139), .A2(n882), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G103), .A2(n524), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U987 ( .A1(n886), .A2(G115), .ZN(n887) );
  XOR2_X1 U988 ( .A(KEYINPUT115), .B(n887), .Z(n890) );
  NAND2_X1 U989 ( .A1(n888), .A2(G127), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n942) );
  XNOR2_X1 U993 ( .A(n894), .B(n942), .ZN(n895) );
  XOR2_X1 U994 ( .A(n896), .B(n895), .Z(n899) );
  XOR2_X1 U995 ( .A(n897), .B(G162), .Z(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U998 ( .A(n903), .B(n902), .Z(n904) );
  NOR2_X1 U999 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT116), .B(n905), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G171), .B(n988), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1003 ( .A(G286), .B(n908), .Z(n909) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1005 ( .A(KEYINPUT110), .B(G2446), .Z(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT111), .B(G2451), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1008 ( .A(KEYINPUT112), .B(G2435), .Z(n913) );
  XNOR2_X1 U1009 ( .A(G2438), .B(G2454), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1012 ( .A(G2443), .B(G2427), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n920) );
  XOR2_X1 U1014 ( .A(G1348), .B(G1341), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G2430), .B(n918), .ZN(n919) );
  XOR2_X1 U1016 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1017 ( .A1(G14), .A2(n921), .ZN(n927) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n927), .ZN(G401) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1029 ( .A(KEYINPUT118), .B(n930), .Z(n931) );
  XNOR2_X1 U1030 ( .A(KEYINPUT51), .B(n931), .ZN(n934) );
  XOR2_X1 U1031 ( .A(G160), .B(G2084), .Z(n932) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n932), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n951) );
  INV_X1 U1034 ( .A(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n949) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G2072), .B(n942), .Z(n944) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT50), .B(n945), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n952), .ZN(n953) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n976), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n954), .A2(G29), .ZN(n1036) );
  XNOR2_X1 U1049 ( .A(KEYINPUT119), .B(G2090), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(G35), .ZN(n974) );
  XNOR2_X1 U1051 ( .A(G2084), .B(G34), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT54), .ZN(n972) );
  XOR2_X1 U1053 ( .A(G2067), .B(G26), .Z(n958) );
  XOR2_X1 U1054 ( .A(G1991), .B(G25), .Z(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n969) );
  XNOR2_X1 U1056 ( .A(G27), .B(n959), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(n960), .B(KEYINPUT121), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G32), .B(n961), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n962), .A2(G28), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT120), .B(G2072), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(G33), .B(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(KEYINPUT53), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1069 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n979), .ZN(n1034) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1007) );
  XNOR2_X1 U1073 ( .A(G168), .B(G1966), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT57), .ZN(n1005) );
  XNOR2_X1 U1076 ( .A(G1956), .B(G299), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(G1961), .B(KEYINPUT123), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n985), .B(G301), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n991) );
  XOR2_X1 U1081 ( .A(G1348), .B(n988), .Z(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n999) );
  XOR2_X1 U1084 ( .A(n992), .B(KEYINPUT124), .Z(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1086 ( .A(G1971), .B(G303), .Z(n995) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT126), .B(n1000), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1032) );
  INV_X1 U1095 ( .A(G16), .ZN(n1030) );
  XNOR2_X1 U1096 ( .A(G20), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G6), .B(G1981), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT59), .B(G1348), .Z(n1013) );
  XNOR2_X1 U1102 ( .A(G4), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G1961), .B(G5), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G1966), .B(G21), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(G1986), .B(G24), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G1971), .B(G22), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1112 ( .A(G1976), .B(G23), .Z(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1121 ( .A(n1037), .B(KEYINPUT127), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1038), .ZN(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

