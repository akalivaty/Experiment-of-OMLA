//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n562, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n463), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(new_n469), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(KEYINPUT67), .B(G2105), .Z(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n473), .A2(new_n480), .A3(new_n482), .ZN(G160));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n478), .C2(G112), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n478), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n475), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n470), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n478), .A2(new_n493), .A3(KEYINPUT4), .A4(G138), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G102), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n493), .A2(new_n495), .B1(new_n498), .B2(G2104), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n511), .B1(new_n505), .B2(new_n506), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(G88), .B1(G50), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n515), .A3(G62), .ZN(new_n516));
  INV_X1    g091(.A(G75), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(new_n511), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n515), .B1(new_n508), .B2(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(G651), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n522), .B(G651), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n514), .B1(new_n521), .B2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(new_n510), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT72), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(G651), .A3(new_n534), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT73), .B(G52), .Z(new_n536));
  AOI22_X1  g111(.A1(new_n510), .A2(G90), .B1(new_n512), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT74), .ZN(G171));
  NAND2_X1  g114(.A1(new_n512), .A2(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n509), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n504), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT75), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n555), .A2(KEYINPUT76), .A3(new_n504), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n510), .A2(G91), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT76), .B1(new_n555), .B2(new_n504), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n554), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  NAND2_X1  g136(.A1(new_n521), .A2(new_n523), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n513), .ZN(G303));
  NAND2_X1  g138(.A1(new_n510), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n512), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(new_n512), .A2(G48), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n508), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n510), .A2(G86), .B1(new_n574), .B2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(G72), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G60), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n504), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(new_n580), .B2(new_n579), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n510), .A2(G85), .B1(G47), .B2(new_n512), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n510), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n572), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(G868), .B2(new_n592), .ZN(G284));
  OAI21_X1  g168(.A(new_n585), .B1(G868), .B2(new_n592), .ZN(G321));
  MUX2_X1   g169(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g170(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g171(.A(KEYINPUT79), .B(G559), .Z(new_n597));
  OAI21_X1  g172(.A(new_n592), .B1(G860), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g174(.A1(new_n592), .A2(new_n597), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n487), .A2(G2104), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT13), .Z(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  OAI221_X1 g187(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n478), .C2(G111), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n485), .A2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n487), .A2(G135), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2096), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(G156));
  XOR2_X1   g193(.A(KEYINPUT15), .B(G2435), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2427), .ZN(new_n621));
  INV_X1    g196(.A(G2430), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n625), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT82), .ZN(new_n633));
  INV_X1    g208(.A(G14), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n630), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT83), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT86), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n643), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n639), .A2(new_n640), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n652));
  OAI221_X1 g227(.A(new_n641), .B1(new_n648), .B2(new_n649), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n610), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n670), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G26), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT28), .Z(new_n679));
  NOR2_X1   g254(.A1(G104), .A2(G2105), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT93), .Z(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(G2104), .C1(G116), .C2(new_n478), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n485), .A2(G128), .B1(new_n487), .B2(G140), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n679), .B1(new_n684), .B2(G29), .ZN(new_n685));
  INV_X1    g260(.A(G2067), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(G4), .A2(G16), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n592), .B2(G16), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n687), .B1(new_n689), .B2(G1348), .ZN(new_n690));
  NOR2_X1   g265(.A1(G16), .A2(G19), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n545), .B2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT92), .B(G1341), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n690), .B(new_n694), .C1(G1348), .C2(new_n689), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT94), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT31), .B(G11), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT30), .B(G28), .Z(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n616), .A2(G29), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g276(.A1(G164), .A2(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G27), .B2(G29), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT101), .B(G2078), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n699), .B(new_n701), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G29), .A2(G35), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G162), .B2(G29), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT29), .Z(new_n709));
  INV_X1    g284(.A(G2090), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n703), .A2(new_n705), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n677), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n485), .A2(G129), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT96), .Z(new_n715));
  AND3_X1   g290(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n716), .B(new_n719), .C1(G141), .C2(new_n487), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n713), .B1(new_n722), .B2(new_n677), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n712), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n727), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1966), .Z(new_n730));
  NAND4_X1  g305(.A1(new_n706), .A2(new_n711), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n709), .A2(new_n710), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT102), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT98), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n723), .A2(new_n725), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n677), .A2(G33), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  NAND2_X1  g312(.A1(G103), .A2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n479), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n478), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n739), .A2(new_n740), .B1(new_n487), .B2(G139), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n493), .A2(G127), .ZN(new_n742));
  AND2_X1   g317(.A1(G115), .A2(G2104), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n479), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n736), .B1(new_n745), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  NAND2_X1  g324(.A1(G160), .A2(G29), .ZN(new_n750));
  AND2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NOR2_X1   g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n677), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(G2084), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n746), .A2(new_n747), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n735), .A2(new_n749), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n731), .B(new_n733), .C1(new_n734), .C2(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n734), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n727), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT23), .Z(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G299), .B2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(G2084), .B1(new_n750), .B2(new_n753), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT100), .Z(new_n765));
  NOR2_X1   g340(.A1(G5), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G171), .B2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(G1961), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n763), .B(new_n768), .C1(G1961), .C2(new_n767), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n696), .A2(new_n757), .A3(new_n758), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n771));
  MUX2_X1   g346(.A(G6), .B(G305), .S(G16), .Z(new_n772));
  XOR2_X1   g347(.A(KEYINPUT32), .B(G1981), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G166), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G16), .B2(G22), .ZN(new_n776));
  INV_X1    g351(.A(G1971), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n727), .A2(G23), .ZN(new_n780));
  INV_X1    g355(.A(G288), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n727), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n774), .A2(new_n778), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT34), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n771), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n787), .A2(KEYINPUT90), .A3(KEYINPUT34), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G290), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G16), .B2(G24), .ZN(new_n796));
  INV_X1    g371(.A(G1986), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR2_X1   g374(.A1(G25), .A2(G29), .ZN(new_n800));
  OAI221_X1 g375(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n478), .C2(G107), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n485), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n487), .A2(G131), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n800), .B1(new_n805), .B2(G29), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n798), .A2(new_n799), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n789), .B2(new_n790), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT91), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n793), .B(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n770), .B1(new_n815), .B2(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(new_n770), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(G150));
  NAND2_X1  g395(.A1(new_n592), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT103), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n510), .A2(G93), .B1(G55), .B2(new_n512), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n504), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n544), .B2(new_n542), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n545), .B(new_n823), .C1(new_n504), .C2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT38), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n822), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT104), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n825), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n721), .B(new_n745), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n684), .B(G164), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n608), .B(new_n804), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n485), .A2(G130), .B1(new_n487), .B2(G142), .ZN(new_n842));
  OAI221_X1 g417(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n478), .C2(G118), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(new_n845), .ZN(new_n847));
  XNOR2_X1  g422(.A(G160), .B(G162), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n616), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT106), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n850), .A2(KEYINPUT106), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n846), .A2(new_n847), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(KEYINPUT105), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n846), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n847), .A2(KEYINPUT105), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n850), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g436(.A1(new_n825), .A2(G868), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n602), .B(new_n828), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n587), .A2(new_n591), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(G299), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(G299), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT107), .B1(new_n867), .B2(KEYINPUT41), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n865), .A2(new_n869), .A3(new_n870), .A4(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(KEYINPUT41), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n867), .B2(new_n863), .ZN(new_n875));
  XNOR2_X1  g450(.A(G166), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(new_n781), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT108), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n876), .A2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n875), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n862), .B1(new_n883), .B2(G868), .ZN(G295));
  AOI21_X1  g459(.A(new_n862), .B1(new_n883), .B2(G868), .ZN(G331));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n886));
  INV_X1    g461(.A(new_n872), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n867), .A2(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(G301), .A2(G286), .ZN(new_n889));
  INV_X1    g464(.A(new_n828), .ZN(new_n890));
  NAND2_X1  g465(.A1(G171), .A2(G168), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n887), .A2(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n865), .A2(new_n866), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n892), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n898), .A3(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n881), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n896), .A2(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n873), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n881), .A3(new_n901), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n854), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n901), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n880), .A3(new_n879), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n854), .A4(new_n906), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n886), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n903), .B2(new_n907), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n910), .A2(KEYINPUT43), .A3(new_n854), .A4(new_n906), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n913), .A2(new_n916), .ZN(G397));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n500), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n473), .A2(G40), .A3(new_n480), .A4(new_n482), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT46), .Z(new_n926));
  INV_X1    g501(.A(new_n923), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n684), .B(new_n686), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n722), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT47), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n794), .A2(new_n797), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT110), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(new_n927), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(KEYINPUT48), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(KEYINPUT48), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n722), .A2(new_n924), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n721), .A2(G1996), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n937), .A2(new_n928), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n805), .A2(new_n807), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n805), .A2(new_n807), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI211_X1 g517(.A(new_n935), .B(new_n936), .C1(new_n923), .C2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n939), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n944), .A2(new_n941), .B1(G2067), .B2(new_n684), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n931), .B(new_n943), .C1(new_n923), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT63), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n918), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND4_X1   g525(.A1(G40), .A2(new_n473), .A3(new_n480), .A4(new_n482), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n500), .A2(KEYINPUT111), .A3(KEYINPUT45), .A4(new_n918), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n950), .A2(new_n921), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n500), .B2(new_n918), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n922), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n950), .A4(new_n952), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n777), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n500), .A2(new_n918), .A3(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n960), .A2(new_n951), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n710), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n959), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(G8), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  NOR3_X1   g547(.A1(G166), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  INV_X1    g551(.A(G1981), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n570), .A2(new_n977), .A3(new_n575), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n977), .B1(new_n570), .B2(new_n575), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n980), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT49), .A3(new_n978), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n922), .A2(new_n919), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT116), .B(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(G288), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n781), .B2(G1976), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n987), .B(new_n990), .C1(new_n989), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n985), .ZN(new_n994));
  INV_X1    g569(.A(G2084), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n960), .A2(new_n951), .A3(new_n995), .A4(new_n962), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1966), .B1(new_n956), .B2(new_n948), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n993), .A2(G286), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n947), .B1(new_n975), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT115), .B1(new_n970), .B2(new_n973), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n971), .B1(G166), .B2(new_n972), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n966), .A2(G8), .A3(new_n1007), .A4(new_n968), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n999), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n500), .A2(new_n1010), .A3(new_n918), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n961), .B1(new_n500), .B2(new_n918), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n922), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n710), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n985), .B1(new_n959), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n974), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n993), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n986), .B(KEYINPUT117), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n987), .A2(new_n988), .A3(new_n781), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n978), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1001), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G168), .A2(new_n985), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n999), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT123), .B1(new_n997), .B2(new_n998), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n921), .A2(new_n951), .A3(new_n948), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1028), .B(new_n996), .C1(new_n1029), .C2(G1966), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(new_n1025), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(new_n1024), .A3(new_n1030), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT51), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1026), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n954), .A2(new_n958), .ZN(new_n1036));
  INV_X1    g611(.A(G2078), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n922), .B1(KEYINPUT50), .B2(new_n919), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1961), .B1(new_n1040), .B2(new_n962), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1037), .A2(KEYINPUT53), .ZN(new_n1042));
  AND4_X1   g617(.A1(new_n921), .A2(new_n951), .A3(new_n948), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n956), .A2(new_n948), .A3(new_n1042), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1045), .B(KEYINPUT124), .C1(new_n963), .C2(G1961), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G171), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n477), .B(KEYINPUT125), .Z(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n478), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n473), .A2(new_n482), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(G40), .ZN(new_n1052));
  NOR4_X1   g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n955), .A4(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n950), .A2(new_n952), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1041), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G2078), .B1(new_n954), .B2(new_n958), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1055), .B(G301), .C1(new_n1056), .C2(KEYINPUT53), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT54), .B1(new_n1048), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1035), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G301), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n1056), .B2(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(G301), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT54), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n959), .A2(new_n1014), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n994), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n993), .B1(new_n1065), .B2(new_n974), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT126), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(new_n1008), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1066), .B2(new_n1008), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1059), .B(new_n1063), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n984), .B2(new_n686), .ZN(new_n1072));
  NOR4_X1   g647(.A1(new_n922), .A2(new_n919), .A3(KEYINPUT120), .A4(G2067), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1040), .A2(new_n962), .ZN(new_n1075));
  INV_X1    g650(.A(G1348), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n864), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT118), .B1(new_n1013), .B2(G1956), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT9), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n512), .B2(G53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(G299), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1080), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n554), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT56), .B(G2072), .Z(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n956), .A2(new_n950), .A3(new_n952), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n500), .A2(new_n1010), .A3(new_n918), .ZN(new_n1095));
  NAND3_X1  g670(.A1(G160), .A2(G40), .A3(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1094), .B(new_n762), .C1(new_n1096), .C2(new_n1012), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1079), .A2(new_n1090), .A3(new_n1093), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1078), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1079), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1090), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1098), .A2(KEYINPUT121), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1098), .A2(KEYINPUT121), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT122), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1105), .B(new_n1110), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n592), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1078), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n953), .A2(G1996), .B1(new_n984), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n545), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(new_n545), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n864), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT61), .B1(new_n1102), .B2(new_n1098), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1103), .B1(new_n1112), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1022), .B1(new_n1070), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1048), .B1(new_n1035), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(KEYINPUT127), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1035), .A2(new_n1129), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1128), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n942), .B1(G1986), .B2(G290), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n927), .B1(new_n1138), .B2(new_n933), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n946), .B1(new_n1137), .B2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g715(.A1(G229), .A2(new_n461), .ZN(new_n1142));
  NAND3_X1  g716(.A1(new_n656), .A2(new_n636), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g717(.A(new_n1143), .B1(new_n859), .B2(new_n855), .ZN(new_n1144));
  AND3_X1   g718(.A1(new_n1144), .A2(new_n914), .A3(new_n915), .ZN(G308));
  NAND3_X1  g719(.A1(new_n1144), .A2(new_n914), .A3(new_n915), .ZN(G225));
endmodule


