//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT25), .B1(new_n208), .B2(KEYINPUT66), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  AOI21_X1  g010(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n212), .A2(KEYINPUT65), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(new_n215), .C1(KEYINPUT65), .C2(new_n212), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n209), .B(new_n216), .C1(KEYINPUT66), .C2(new_n208), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT27), .B(G183gat), .Z(new_n218));
  OAI21_X1  g017(.A(KEYINPUT28), .B1(new_n218), .B2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n213), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT27), .B1(new_n213), .B2(KEYINPUT69), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n219), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT70), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n207), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n207), .B(KEYINPUT67), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n210), .B1(new_n212), .B2(KEYINPUT68), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n212), .A2(new_n210), .A3(KEYINPUT68), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n206), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n225), .A2(new_n229), .B1(new_n234), .B2(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n236), .A2(G226gat), .A3(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n236), .A2(new_n238), .B1(G226gat), .B2(G233gat), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G197gat), .B(G204gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT74), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n242), .A2(new_n243), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n248), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n240), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n237), .A2(new_n239), .ZN(new_n253));
  INV_X1    g052(.A(new_n251), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G64gat), .B(G92gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT76), .ZN(new_n258));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  OR2_X1    g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n260), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(KEYINPUT30), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT30), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n256), .A2(new_n264), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT1), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G141gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G148gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT78), .B(G148gat), .Z(new_n279));
  OAI211_X1 g078(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n274), .ZN(new_n280));
  XNOR2_X1  g079(.A(G155gat), .B(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT79), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(G155gat), .B2(G162gat), .ZN(new_n284));
  XOR2_X1   g083(.A(G155gat), .B(G162gat), .Z(new_n285));
  INV_X1    g084(.A(KEYINPUT79), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n280), .A2(new_n287), .A3(KEYINPUT80), .A4(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G148gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G141gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n281), .B1(new_n295), .B2(new_n283), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n273), .B1(new_n299), .B2(KEYINPUT81), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n296), .B1(new_n290), .B2(new_n291), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI211_X1 g103(.A(KEYINPUT3), .B(new_n296), .C1(new_n290), .C2(new_n291), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n268), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT5), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n273), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT4), .ZN(new_n311));
  AOI211_X1 g110(.A(new_n296), .B(new_n272), .C1(new_n290), .C2(new_n291), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(KEYINPUT84), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT89), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n303), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT81), .B1(new_n299), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n272), .B1(new_n304), .B2(new_n301), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n267), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n326), .A3(KEYINPUT4), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT82), .B1(new_n312), .B2(new_n313), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n310), .A2(KEYINPUT4), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n325), .A2(KEYINPUT83), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n312), .A2(KEYINPUT82), .A3(new_n313), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n326), .B1(new_n310), .B2(KEYINPUT4), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(new_n314), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n307), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n302), .A2(new_n273), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n312), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT5), .B1(new_n339), .B2(new_n267), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n320), .B(new_n321), .C1(new_n337), .C2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT83), .B1(new_n325), .B2(new_n330), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n307), .A2(new_n335), .A3(new_n332), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT89), .B1(new_n344), .B2(new_n319), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  INV_X1    g145(.A(G85gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G57gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n344), .A2(new_n319), .ZN(new_n352));
  INV_X1    g151(.A(new_n350), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT6), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(KEYINPUT6), .B(new_n350), .C1(new_n344), .C2(new_n319), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n202), .B(new_n266), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n251), .B1(new_n322), .B2(new_n238), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n246), .B2(new_n250), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n250), .B2(new_n246), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n302), .B1(new_n303), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n364), .B(KEYINPUT85), .Z(new_n365));
  NAND2_X1  g164(.A1(new_n251), .A2(new_n238), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n366), .A2(KEYINPUT86), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n303), .B1(new_n366), .B2(KEYINPUT86), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n298), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n359), .A2(new_n364), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n363), .A2(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(G22gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT31), .B(G50gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(new_n375), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(KEYINPUT35), .ZN(new_n379));
  XNOR2_X1  g178(.A(G15gat), .B(G43gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g181(.A(G227gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n236), .A2(new_n272), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n217), .A2(new_n273), .A3(new_n235), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n382), .B1(new_n389), .B2(KEYINPUT33), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT32), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n392), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(new_n386), .A3(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT34), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT34), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n387), .A2(new_n398), .A3(new_n386), .A4(new_n388), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(new_n394), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT91), .B1(new_n401), .B2(new_n403), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n379), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n357), .B1(new_n351), .B2(new_n354), .ZN(new_n410));
  INV_X1    g209(.A(new_n266), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT90), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n358), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n350), .B1(new_n344), .B2(new_n319), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n354), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n415), .B2(new_n356), .ZN(new_n416));
  INV_X1    g215(.A(new_n378), .ZN(new_n417));
  INV_X1    g216(.A(new_n394), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n390), .A2(new_n392), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n397), .B2(new_n399), .ZN(new_n422));
  OAI22_X1  g221(.A1(new_n418), .A2(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT72), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n395), .B(new_n425), .C1(new_n422), .C2(new_n420), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n417), .A2(new_n424), .A3(new_n426), .A4(new_n403), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n256), .A2(KEYINPUT37), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n252), .A2(new_n431), .A3(new_n255), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n260), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT38), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n262), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n434), .B2(new_n433), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n378), .B1(new_n436), .B2(new_n410), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n316), .B(new_n317), .C1(new_n323), .C2(new_n324), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n268), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n339), .B2(new_n267), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n440), .A3(new_n268), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n443), .A2(new_n444), .A3(new_n353), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n443), .B2(new_n353), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n447), .A2(KEYINPUT88), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT88), .B1(new_n447), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n411), .B(new_n351), .C1(new_n448), .C2(new_n447), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n437), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  INV_X1    g253(.A(new_n403), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n402), .B1(new_n393), .B2(new_n394), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT36), .A4(new_n403), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n404), .A2(KEYINPUT73), .A3(new_n454), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n415), .A2(new_n356), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n266), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(new_n378), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n413), .A2(new_n429), .B1(new_n453), .B2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G15gat), .B(G22gat), .Z(new_n467));
  INV_X1    g266(.A(G1gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n468), .A2(KEYINPUT16), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n469), .B(KEYINPUT98), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G8gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(G57gat), .B(G64gat), .Z(new_n474));
  INV_X1    g273(.A(KEYINPUT9), .ZN(new_n475));
  INV_X1    g274(.A(G71gat), .ZN(new_n476));
  INV_X1    g275(.A(G78gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT21), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n482), .A2(KEYINPUT21), .A3(new_n481), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n473), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n473), .B2(new_n483), .ZN(new_n486));
  XNOR2_X1  g285(.A(G127gat), .B(G155gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G231gat), .A2(G233gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(new_n213), .ZN(new_n492));
  INV_X1    g291(.A(G211gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n490), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT15), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n499), .B2(new_n498), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n502));
  INV_X1    g301(.A(G29gat), .ZN(new_n503));
  INV_X1    g302(.A(G36gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT97), .B(KEYINPUT15), .ZN(new_n508));
  OAI221_X1 g307(.A(new_n507), .B1(new_n503), .B2(new_n504), .C1(new_n498), .C2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n507), .A2(KEYINPUT95), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n501), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n501), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT17), .B(new_n510), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  AND2_X1   g320(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n522));
  NOR2_X1   g321(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n523));
  INV_X1    g322(.A(G92gat), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n522), .A2(new_n523), .B1(new_n347), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT102), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  AOI22_X1  g331(.A1(KEYINPUT8), .A2(new_n532), .B1(new_n347), .B2(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G99gat), .B(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n525), .A2(new_n531), .A3(new_n535), .A4(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT103), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n521), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n541), .ZN(new_n544));
  INV_X1    g343(.A(G232gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n384), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT104), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT104), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  AOI211_X1 g349(.A(new_n549), .B(new_n550), .C1(new_n518), .C2(new_n541), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n543), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT101), .ZN(new_n556));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n553), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(new_n543), .C1(new_n548), .C2(new_n551), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n558), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n497), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n466), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n473), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n518), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n521), .A2(new_n473), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n501), .A2(new_n514), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT96), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n501), .A2(new_n514), .A3(new_n515), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT17), .B1(new_n574), .B2(new_n510), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n567), .B(new_n569), .C1(new_n570), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n520), .A2(new_n473), .A3(new_n521), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n567), .A4(new_n569), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n567), .B(KEYINPUT13), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n569), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n518), .A2(new_n568), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n578), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n586), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n578), .A2(new_n593), .A3(new_n580), .A4(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n541), .A2(KEYINPUT10), .A3(new_n482), .A4(new_n481), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT105), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n539), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n481), .A2(new_n482), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n537), .A2(KEYINPUT105), .A3(new_n538), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n539), .A2(new_n600), .A3(new_n482), .A4(new_n481), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT106), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT106), .ZN(new_n609));
  AOI211_X1 g408(.A(new_n609), .B(KEYINPUT10), .C1(new_n604), .C2(new_n605), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n599), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n604), .A2(new_n614), .A3(new_n605), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n613), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n598), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n566), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n463), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n468), .ZN(G1324gat));
  NOR2_X1   g426(.A1(new_n625), .A2(new_n266), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n472), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT16), .B(G8gat), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n633), .B2(KEYINPUT42), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(KEYINPUT42), .B2(new_n633), .ZN(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n625), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n406), .A2(new_n407), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n636), .B2(new_n640), .ZN(G1326gat));
  NAND3_X1  g440(.A1(new_n566), .A2(new_n624), .A3(new_n378), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT108), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT43), .B(G22gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  NOR2_X1   g444(.A1(new_n466), .A2(new_n564), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n497), .A2(new_n598), .A3(new_n623), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n648), .A2(G29gat), .A3(new_n463), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT45), .Z(new_n650));
  NOR2_X1   g449(.A1(new_n410), .A2(new_n411), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n408), .B1(new_n651), .B2(new_n202), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n652), .A2(new_n412), .B1(KEYINPUT35), .B2(new_n428), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n637), .B1(new_n416), .B2(new_n417), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n452), .A2(new_n451), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n437), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n563), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n497), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(KEYINPUT44), .B(new_n563), .C1(new_n653), .C2(new_n656), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n624), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(G29gat), .B1(new_n661), .B2(new_n463), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n650), .A2(new_n662), .ZN(G1328gat));
  NOR3_X1   g462(.A1(new_n648), .A2(G36gat), .A3(new_n266), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT46), .ZN(new_n665));
  OAI21_X1  g464(.A(G36gat), .B1(new_n661), .B2(new_n266), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(G1329gat));
  NAND2_X1  g466(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n668));
  INV_X1    g467(.A(G43gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n648), .B2(new_n639), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n462), .A2(G43gat), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n668), .B(new_n670), .C1(new_n661), .C2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(G1330gat));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n417), .B1(new_n648), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n646), .A2(KEYINPUT110), .A3(new_n647), .ZN(new_n677));
  AOI21_X1  g476(.A(G50gat), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n378), .A2(G50gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n679), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n678), .A2(new_n680), .A3(KEYINPUT48), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT48), .B1(new_n678), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1331gat));
  INV_X1    g482(.A(new_n623), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n597), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n566), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n463), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n266), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  AND2_X1   g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n689), .B2(new_n690), .ZN(G1333gat));
  OAI21_X1  g492(.A(new_n476), .B1(new_n686), .B2(new_n639), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n462), .A2(G71gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n686), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1334gat));
  NOR2_X1   g497(.A1(new_n686), .A2(new_n417), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(new_n477), .ZN(G1335gat));
  NOR2_X1   g499(.A1(new_n497), .A2(new_n597), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n646), .A2(KEYINPUT51), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n657), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n463), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n706), .A2(new_n347), .A3(new_n707), .A4(new_n623), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n658), .B1(new_n466), .B2(new_n564), .ZN(new_n709));
  INV_X1    g508(.A(new_n497), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n660), .A3(new_n710), .A4(new_n685), .ZN(new_n711));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711), .B2(new_n463), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(G1336gat));
  NAND4_X1  g512(.A1(new_n706), .A2(new_n524), .A3(new_n623), .A4(new_n411), .ZN(new_n714));
  OAI21_X1  g513(.A(G92gat), .B1(new_n711), .B2(new_n266), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n711), .B2(new_n637), .ZN(new_n718));
  INV_X1    g517(.A(new_n706), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n639), .A2(G99gat), .A3(new_n684), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT112), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n719), .B2(new_n721), .ZN(G1338gat));
  OAI21_X1  g521(.A(G106gat), .B1(new_n711), .B2(new_n417), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT113), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n725), .B(G106gat), .C1(new_n711), .C2(new_n417), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n417), .A2(G106gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n706), .A2(KEYINPUT114), .A3(new_n623), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n724), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT53), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n623), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(KEYINPUT114), .A2(KEYINPUT53), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n731), .B(new_n732), .C1(new_n723), .C2(KEYINPUT53), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(G1339gat));
  NAND4_X1  g533(.A1(new_n497), .A2(new_n598), .A3(new_n684), .A4(new_n564), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n614), .B(new_n599), .C1(new_n608), .C2(new_n610), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n613), .A2(KEYINPUT54), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT54), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n611), .A2(new_n739), .A3(new_n612), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n738), .A2(KEYINPUT55), .A3(new_n619), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n622), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT115), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n622), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(new_n619), .A3(new_n740), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n567), .B1(new_n579), .B2(new_n569), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n583), .A2(new_n584), .A3(new_n582), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n591), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n596), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n561), .A2(new_n752), .A3(new_n562), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n743), .A2(new_n745), .A3(new_n748), .A4(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n742), .A2(KEYINPUT115), .B1(new_n747), .B2(new_n746), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(KEYINPUT116), .A3(new_n745), .A4(new_n753), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n597), .A3(new_n745), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n623), .A2(new_n596), .A3(new_n751), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(new_n563), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n736), .B1(new_n763), .B2(new_n710), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n378), .A3(new_n639), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n463), .A2(new_n411), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G113gat), .B1(new_n767), .B2(new_n598), .ZN(new_n768));
  INV_X1    g567(.A(new_n764), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n427), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n766), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n598), .A2(G113gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(G1340gat));
  OAI21_X1  g572(.A(G120gat), .B1(new_n767), .B2(new_n684), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n684), .A2(G120gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n771), .B2(new_n775), .ZN(G1341gat));
  INV_X1    g575(.A(G127gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n767), .A2(new_n777), .A3(new_n710), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n770), .A2(new_n497), .A3(new_n766), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(G1342gat));
  OR2_X1    g579(.A1(new_n564), .A2(G134gat), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n771), .A2(KEYINPUT56), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n563), .A3(new_n766), .A4(new_n769), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G134gat), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT56), .B1(new_n771), .B2(new_n781), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(G1343gat));
  INV_X1    g585(.A(KEYINPUT121), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n417), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n748), .A2(new_n597), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n761), .B1(new_n790), .B2(new_n742), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n564), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n497), .B1(new_n759), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n735), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g594(.A(KEYINPUT118), .B(new_n497), .C1(new_n759), .C2(new_n792), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT119), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(new_n789), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n756), .A2(new_n758), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n563), .B1(new_n760), .B2(new_n761), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n710), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n417), .B1(new_n803), .B2(new_n735), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT117), .B1(new_n804), .B2(KEYINPUT57), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n806), .B(new_n788), .C1(new_n764), .C2(new_n417), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n798), .A2(new_n800), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n462), .A2(new_n463), .A3(new_n411), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n597), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G141gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n804), .A2(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n597), .A2(new_n274), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n787), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g616(.A(KEYINPUT121), .B(new_n815), .C1(new_n810), .C2(G141gat), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n813), .A2(new_n814), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(G141gat), .B2(new_n810), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n817), .A2(new_n818), .B1(new_n812), .B2(new_n822), .ZN(G1344gat));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n824), .B(new_n279), .C1(new_n825), .C2(new_n684), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT57), .B1(new_n764), .B2(new_n417), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n735), .B(KEYINPUT122), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n497), .B1(new_n792), .B2(new_n754), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n788), .B(new_n378), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n623), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n293), .B1(new_n832), .B2(new_n809), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n826), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n684), .A2(new_n279), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n813), .B2(new_n835), .ZN(G1345gat));
  NAND4_X1  g635(.A1(new_n808), .A2(G155gat), .A3(new_n497), .A4(new_n809), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n804), .A2(new_n497), .A3(new_n809), .ZN(new_n838));
  AOI21_X1  g637(.A(G155gat), .B1(new_n838), .B2(KEYINPUT123), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(KEYINPUT123), .B2(new_n838), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n837), .A2(new_n840), .ZN(G1346gat));
  NAND2_X1  g640(.A1(new_n563), .A2(G162gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n813), .A2(new_n564), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n825), .A2(new_n842), .B1(G162gat), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT124), .ZN(G1347gat));
  NOR2_X1   g644(.A1(new_n707), .A2(new_n266), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n765), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G169gat), .B1(new_n847), .B2(new_n598), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n770), .A2(new_n846), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n597), .A2(new_n203), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1348gat));
  NOR3_X1   g650(.A1(new_n847), .A2(new_n204), .A3(new_n684), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n770), .A2(new_n623), .A3(new_n846), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n204), .B2(new_n853), .ZN(G1349gat));
  OAI21_X1  g653(.A(G183gat), .B1(new_n847), .B2(new_n710), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n710), .A2(new_n218), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g657(.A1(new_n765), .A2(new_n563), .A3(new_n846), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(G190gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(G190gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n563), .A2(new_n214), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n861), .A2(new_n862), .B1(new_n849), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT125), .ZN(G1351gat));
  NOR3_X1   g664(.A1(new_n707), .A2(new_n462), .A3(new_n266), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n831), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G197gat), .B1(new_n867), .B2(new_n598), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n804), .A2(new_n866), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n598), .A2(G197gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(G1352gat));
  NAND2_X1  g670(.A1(new_n832), .A2(new_n866), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G204gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n869), .A2(G204gat), .A3(new_n684), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT62), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1353gat));
  OAI21_X1  g675(.A(G211gat), .B1(new_n867), .B2(new_n710), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT63), .B(G211gat), .C1(new_n867), .C2(new_n710), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n497), .A2(new_n493), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n882), .A2(new_n883), .B1(new_n869), .B2(new_n884), .ZN(G1354gat));
  NAND2_X1  g684(.A1(new_n563), .A2(G218gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n564), .ZN(new_n887));
  OAI22_X1  g686(.A1(new_n867), .A2(new_n886), .B1(G218gat), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT127), .Z(G1355gat));
endmodule


