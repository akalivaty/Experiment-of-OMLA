

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786;

  AND2_X1 U381 ( .A1(n409), .A2(n406), .ZN(n373) );
  INV_X1 U382 ( .A(n617), .ZN(n702) );
  XNOR2_X2 U383 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n420) );
  NAND2_X2 U384 ( .A1(n373), .A2(n377), .ZN(n400) );
  AND2_X2 U385 ( .A1(n403), .A2(n379), .ZN(n401) );
  OR2_X2 U386 ( .A1(n404), .A2(n402), .ZN(n379) );
  NOR2_X2 U387 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X2 U388 ( .A(n477), .B(n421), .ZN(n458) );
  NOR2_X1 U389 ( .A1(n611), .A2(n708), .ZN(n612) );
  INV_X2 U390 ( .A(G953), .ZN(n781) );
  XNOR2_X1 U391 ( .A(n514), .B(n513), .ZN(n785) );
  XNOR2_X1 U392 ( .A(n534), .B(KEYINPUT78), .ZN(n674) );
  INV_X1 U393 ( .A(n602), .ZN(n365) );
  NAND2_X1 U394 ( .A1(n755), .A2(n751), .ZN(n718) );
  AND2_X1 U395 ( .A1(n541), .A2(n540), .ZN(n714) );
  AND2_X1 U396 ( .A1(n364), .A2(n363), .ZN(n362) );
  INV_X1 U397 ( .A(KEYINPUT16), .ZN(n358) );
  INV_X1 U398 ( .A(KEYINPUT102), .ZN(n372) );
  NOR2_X1 U399 ( .A1(n693), .A2(n641), .ZN(n695) );
  INV_X1 U400 ( .A(n746), .ZN(n368) );
  AND2_X1 U401 ( .A1(n596), .A2(n593), .ZN(n595) );
  NAND2_X1 U402 ( .A1(n365), .A2(n588), .ZN(n590) );
  OR2_X1 U403 ( .A1(n729), .A2(n533), .ZN(n527) );
  XNOR2_X1 U404 ( .A(n609), .B(n372), .ZN(n370) );
  NOR2_X1 U405 ( .A1(n432), .A2(n518), .ZN(n542) );
  NAND2_X1 U406 ( .A1(n543), .A2(n717), .ZN(n367) );
  NAND2_X2 U407 ( .A1(n362), .A2(n360), .ZN(n543) );
  XNOR2_X1 U408 ( .A(n384), .B(n451), .ZN(n617) );
  XNOR2_X1 U409 ( .A(n497), .B(n496), .ZN(n541) );
  OR2_X1 U410 ( .A1(n664), .A2(G902), .ZN(n384) );
  XNOR2_X1 U411 ( .A(n761), .B(n478), .ZN(n645) );
  OR2_X1 U412 ( .A1(n480), .A2(n629), .ZN(n361) );
  NAND2_X1 U413 ( .A1(n480), .A2(n629), .ZN(n363) );
  XNOR2_X1 U414 ( .A(n503), .B(n420), .ZN(n477) );
  XNOR2_X1 U415 ( .A(G119), .B(G113), .ZN(n416) );
  XNOR2_X1 U416 ( .A(G101), .B(KEYINPUT67), .ZN(n415) );
  XNOR2_X1 U417 ( .A(G146), .B(G125), .ZN(n472) );
  XNOR2_X1 U418 ( .A(G104), .B(G122), .ZN(n485) );
  XNOR2_X1 U419 ( .A(G110), .B(KEYINPUT74), .ZN(n468) );
  XNOR2_X1 U420 ( .A(G116), .B(G107), .ZN(n504) );
  XNOR2_X1 U421 ( .A(n359), .B(n357), .ZN(n470) );
  XNOR2_X1 U422 ( .A(n468), .B(n358), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n485), .B(n504), .ZN(n359) );
  OR2_X1 U424 ( .A1(n645), .A2(n361), .ZN(n360) );
  NAND2_X1 U425 ( .A1(n645), .A2(n480), .ZN(n364) );
  NAND2_X1 U426 ( .A1(n365), .A2(n604), .ZN(n410) );
  NAND2_X1 U427 ( .A1(n365), .A2(n614), .ZN(n743) );
  NOR2_X1 U428 ( .A1(n376), .A2(n366), .ZN(n605) );
  NOR2_X1 U429 ( .A1(n366), .A2(n606), .ZN(n607) );
  NAND2_X1 U430 ( .A1(n369), .A2(n368), .ZN(n366) );
  NAND2_X1 U431 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X2 U432 ( .A(n367), .B(KEYINPUT19), .ZN(n584) );
  INV_X1 U433 ( .A(n786), .ZN(n369) );
  NAND2_X1 U434 ( .A1(n370), .A2(n599), .ZN(n601) );
  NAND2_X2 U435 ( .A1(n371), .A2(n698), .ZN(n609) );
  INV_X1 U436 ( .A(n598), .ZN(n371) );
  AND2_X1 U437 ( .A1(n643), .A2(n642), .ZN(n685) );
  OR2_X2 U438 ( .A1(n712), .A2(n410), .ZN(n409) );
  XNOR2_X1 U439 ( .A(n632), .B(KEYINPUT64), .ZN(n643) );
  AND2_X2 U440 ( .A1(n643), .A2(n642), .ZN(n374) );
  BUF_X1 U441 ( .A(n609), .Z(n375) );
  NAND2_X1 U442 ( .A1(n401), .A2(n400), .ZN(n376) );
  NAND2_X1 U443 ( .A1(n401), .A2(n400), .ZN(n678) );
  XNOR2_X2 U444 ( .A(n774), .B(n466), .ZN(n687) );
  XNOR2_X2 U445 ( .A(n458), .B(n457), .ZN(n774) );
  OR2_X1 U446 ( .A1(n674), .A2(n556), .ZN(n557) );
  OR2_X1 U447 ( .A1(n674), .A2(n539), .ZN(n553) );
  AND2_X1 U448 ( .A1(n553), .A2(n552), .ZN(n559) );
  XNOR2_X1 U449 ( .A(G128), .B(G119), .ZN(n438) );
  XNOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n436) );
  NAND2_X1 U451 ( .A1(n389), .A2(n386), .ZN(n385) );
  AND2_X1 U452 ( .A1(n387), .A2(n629), .ZN(n386) );
  NAND2_X1 U453 ( .A1(n634), .A2(n380), .ZN(n389) );
  NAND2_X1 U454 ( .A1(n388), .A2(n579), .ZN(n387) );
  AND2_X1 U455 ( .A1(n407), .A2(n378), .ZN(n406) );
  INV_X1 U456 ( .A(G101), .ZN(n461) );
  XNOR2_X1 U457 ( .A(G107), .B(G146), .ZN(n462) );
  INV_X1 U458 ( .A(KEYINPUT35), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n524), .B(KEYINPUT103), .ZN(n382) );
  XNOR2_X1 U460 ( .A(n523), .B(n522), .ZN(n383) );
  INV_X1 U461 ( .A(n578), .ZN(n388) );
  NAND2_X1 U462 ( .A1(n394), .A2(n393), .ZN(n392) );
  NOR2_X1 U463 ( .A1(n569), .A2(n570), .ZN(n394) );
  INV_X1 U464 ( .A(KEYINPUT45), .ZN(n626) );
  XNOR2_X1 U465 ( .A(G110), .B(KEYINPUT91), .ZN(n437) );
  XNOR2_X1 U466 ( .A(n445), .B(n444), .ZN(n498) );
  XNOR2_X1 U467 ( .A(G143), .B(G113), .ZN(n483) );
  XNOR2_X1 U468 ( .A(n472), .B(n442), .ZN(n775) );
  INV_X1 U469 ( .A(KEYINPUT66), .ZN(n441) );
  NAND2_X1 U470 ( .A1(n617), .A2(n520), .ZN(n562) );
  INV_X1 U471 ( .A(G902), .ZN(n509) );
  AND2_X1 U472 ( .A1(n698), .A2(n566), .ZN(n544) );
  XNOR2_X1 U473 ( .A(n585), .B(KEYINPUT0), .ZN(n602) );
  XNOR2_X1 U474 ( .A(G116), .B(G146), .ZN(n411) );
  XOR2_X1 U475 ( .A(G137), .B(KEYINPUT5), .Z(n412) );
  NAND2_X1 U476 ( .A1(n634), .A2(n578), .ZN(n780) );
  NAND2_X1 U477 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U478 ( .A1(n719), .A2(n515), .ZN(n517) );
  OR2_X1 U479 ( .A1(n616), .A2(n395), .ZN(n574) );
  NAND2_X1 U480 ( .A1(n398), .A2(n396), .ZN(n395) );
  NOR2_X1 U481 ( .A1(n562), .A2(n397), .ZN(n396) );
  AND2_X1 U482 ( .A1(n382), .A2(n584), .ZN(n381) );
  NAND2_X1 U483 ( .A1(n399), .A2(n540), .ZN(n751) );
  INV_X1 U484 ( .A(n751), .ZN(n398) );
  AND2_X1 U485 ( .A1(n404), .A2(n402), .ZN(n377) );
  NOR2_X1 U486 ( .A1(n541), .A2(n540), .ZN(n378) );
  AND2_X1 U487 ( .A1(n578), .A2(KEYINPUT75), .ZN(n380) );
  XNOR2_X1 U488 ( .A(n511), .B(n510), .ZN(n540) );
  BUF_X1 U489 ( .A(n602), .Z(n611) );
  INV_X1 U490 ( .A(n717), .ZN(n397) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n580) );
  NAND2_X1 U492 ( .A1(n383), .A2(n382), .ZN(n533) );
  NAND2_X1 U493 ( .A1(n381), .A2(n383), .ZN(n534) );
  XNOR2_X1 U494 ( .A(n450), .B(n449), .ZN(n664) );
  NOR2_X1 U495 ( .A1(n390), .A2(n385), .ZN(n391) );
  NOR2_X1 U496 ( .A1(n634), .A2(KEYINPUT75), .ZN(n390) );
  NAND2_X1 U497 ( .A1(n633), .A2(n391), .ZN(n628) );
  XNOR2_X1 U498 ( .A(n532), .B(n531), .ZN(n393) );
  XNOR2_X2 U499 ( .A(n392), .B(n571), .ZN(n634) );
  INV_X1 U500 ( .A(n541), .ZN(n399) );
  NAND2_X1 U501 ( .A1(n405), .A2(KEYINPUT35), .ZN(n403) );
  NAND2_X1 U502 ( .A1(n712), .A2(n408), .ZN(n404) );
  NAND2_X1 U503 ( .A1(n409), .A2(n406), .ZN(n405) );
  NAND2_X1 U504 ( .A1(n611), .A2(n408), .ZN(n407) );
  INV_X1 U505 ( .A(n604), .ZN(n408) );
  XNOR2_X1 U506 ( .A(n627), .B(n626), .ZN(n633) );
  BUF_X1 U507 ( .A(n633), .Z(n765) );
  XNOR2_X1 U508 ( .A(n566), .B(n565), .ZN(n598) );
  INV_X1 U509 ( .A(KEYINPUT75), .ZN(n579) );
  INV_X1 U510 ( .A(n695), .ZN(n642) );
  XNOR2_X1 U511 ( .A(n423), .B(G472), .ZN(n561) );
  BUF_X1 U512 ( .A(n561), .Z(n705) );
  INV_X1 U513 ( .A(KEYINPUT122), .ZN(n668) );
  INV_X1 U514 ( .A(KEYINPUT30), .ZN(n426) );
  XNOR2_X1 U515 ( .A(n412), .B(n411), .ZN(n414) );
  NOR2_X1 U516 ( .A1(G953), .A2(G237), .ZN(n490) );
  NAND2_X1 U517 ( .A1(n490), .A2(G210), .ZN(n413) );
  XNOR2_X1 U518 ( .A(n414), .B(n413), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n416), .B(n415), .ZN(n418) );
  XNOR2_X1 U520 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n418), .B(n417), .ZN(n469) );
  XNOR2_X1 U522 ( .A(n419), .B(n469), .ZN(n422) );
  XNOR2_X2 U523 ( .A(G143), .B(G128), .ZN(n503) );
  XNOR2_X1 U524 ( .A(G134), .B(G131), .ZN(n421) );
  XNOR2_X1 U525 ( .A(n422), .B(n458), .ZN(n680) );
  NAND2_X1 U526 ( .A1(n680), .A2(n509), .ZN(n423) );
  INV_X1 U527 ( .A(G237), .ZN(n424) );
  NAND2_X1 U528 ( .A1(n509), .A2(n424), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n479), .A2(G214), .ZN(n717) );
  AND2_X1 U530 ( .A1(n561), .A2(n717), .ZN(n425) );
  XNOR2_X1 U531 ( .A(n426), .B(n425), .ZN(n432) );
  NAND2_X1 U532 ( .A1(G237), .A2(G234), .ZN(n427) );
  XNOR2_X1 U533 ( .A(n427), .B(KEYINPUT14), .ZN(n697) );
  NOR2_X1 U534 ( .A1(G902), .A2(n781), .ZN(n429) );
  NOR2_X1 U535 ( .A1(G953), .A2(G952), .ZN(n428) );
  NOR2_X1 U536 ( .A1(n429), .A2(n428), .ZN(n430) );
  AND2_X1 U537 ( .A1(n697), .A2(n430), .ZN(n582) );
  NAND2_X1 U538 ( .A1(G953), .A2(G900), .ZN(n431) );
  NAND2_X1 U539 ( .A1(n582), .A2(n431), .ZN(n518) );
  NAND2_X1 U540 ( .A1(n580), .A2(G234), .ZN(n433) );
  XNOR2_X1 U541 ( .A(n433), .B(KEYINPUT92), .ZN(n434) );
  XNOR2_X1 U542 ( .A(n434), .B(KEYINPUT20), .ZN(n452) );
  NAND2_X1 U543 ( .A1(n452), .A2(G217), .ZN(n435) );
  XNOR2_X1 U544 ( .A(n435), .B(KEYINPUT25), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n437), .B(n436), .ZN(n440) );
  XNOR2_X1 U546 ( .A(n438), .B(KEYINPUT81), .ZN(n439) );
  XNOR2_X1 U547 ( .A(n440), .B(n439), .ZN(n443) );
  XNOR2_X1 U548 ( .A(n441), .B(KEYINPUT10), .ZN(n442) );
  XNOR2_X1 U549 ( .A(n443), .B(n775), .ZN(n450) );
  NAND2_X1 U550 ( .A1(G234), .A2(n781), .ZN(n445) );
  INV_X1 U551 ( .A(KEYINPUT8), .ZN(n444) );
  NAND2_X1 U552 ( .A1(n498), .A2(G221), .ZN(n448) );
  XNOR2_X1 U553 ( .A(G137), .B(G140), .ZN(n456) );
  XNOR2_X1 U554 ( .A(KEYINPUT69), .B(KEYINPUT76), .ZN(n446) );
  XNOR2_X1 U555 ( .A(n456), .B(n446), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U557 ( .A1(n452), .A2(G221), .ZN(n454) );
  INV_X1 U558 ( .A(KEYINPUT21), .ZN(n453) );
  XNOR2_X1 U559 ( .A(n454), .B(n453), .ZN(n701) );
  INV_X1 U560 ( .A(KEYINPUT93), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n701), .B(n455), .ZN(n586) );
  AND2_X1 U562 ( .A1(n702), .A2(n586), .ZN(n698) );
  XNOR2_X1 U563 ( .A(n456), .B(KEYINPUT89), .ZN(n457) );
  NAND2_X1 U564 ( .A1(n781), .A2(G227), .ZN(n459) );
  XNOR2_X1 U565 ( .A(n459), .B(KEYINPUT90), .ZN(n460) );
  XNOR2_X1 U566 ( .A(n460), .B(n468), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n461), .B(G104), .ZN(n463) );
  XNOR2_X1 U568 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n465), .B(n464), .ZN(n466) );
  OR2_X2 U570 ( .A1(n687), .A2(G902), .ZN(n467) );
  XNOR2_X2 U571 ( .A(n467), .B(G469), .ZN(n566) );
  NAND2_X1 U572 ( .A1(n542), .A2(n544), .ZN(n481) );
  XNOR2_X1 U573 ( .A(n470), .B(n469), .ZN(n761) );
  XNOR2_X1 U574 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n472), .B(n471), .ZN(n475) );
  NAND2_X1 U576 ( .A1(n781), .A2(G224), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n473), .B(KEYINPUT87), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U580 ( .A(n580), .ZN(n629) );
  AND2_X1 U581 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U582 ( .A(n543), .B(KEYINPUT38), .ZN(n719) );
  OR2_X2 U583 ( .A1(n481), .A2(n719), .ZN(n482) );
  XNOR2_X2 U584 ( .A(n482), .B(KEYINPUT39), .ZN(n573) );
  XOR2_X1 U585 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n484) );
  XNOR2_X1 U586 ( .A(n484), .B(n483), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U588 ( .A(n487), .B(n775), .ZN(n495) );
  XOR2_X1 U589 ( .A(G131), .B(KEYINPUT94), .Z(n489) );
  XNOR2_X1 U590 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U591 ( .A(n489), .B(n488), .ZN(n493) );
  NAND2_X1 U592 ( .A1(n490), .A2(G214), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n491), .B(G140), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U595 ( .A(n495), .B(n494), .ZN(n653) );
  NAND2_X1 U596 ( .A1(n653), .A2(n509), .ZN(n497) );
  XNOR2_X1 U597 ( .A(KEYINPUT13), .B(G475), .ZN(n496) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n500) );
  NAND2_X1 U599 ( .A1(G217), .A2(n498), .ZN(n499) );
  XNOR2_X1 U600 ( .A(n500), .B(n499), .ZN(n508) );
  XOR2_X1 U601 ( .A(G134), .B(KEYINPUT98), .Z(n502) );
  XNOR2_X1 U602 ( .A(G122), .B(KEYINPUT7), .ZN(n501) );
  XNOR2_X1 U603 ( .A(n502), .B(n501), .ZN(n506) );
  XNOR2_X1 U604 ( .A(n503), .B(n504), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U606 ( .A(n508), .B(n507), .ZN(n659) );
  NAND2_X1 U607 ( .A1(n659), .A2(n509), .ZN(n511) );
  XNOR2_X1 U608 ( .A(G478), .B(KEYINPUT99), .ZN(n510) );
  INV_X1 U609 ( .A(n540), .ZN(n535) );
  NAND2_X1 U610 ( .A1(n573), .A2(n398), .ZN(n514) );
  INV_X1 U611 ( .A(KEYINPUT104), .ZN(n512) );
  XNOR2_X1 U612 ( .A(n512), .B(KEYINPUT40), .ZN(n513) );
  INV_X1 U613 ( .A(n785), .ZN(n529) );
  NAND2_X1 U614 ( .A1(n714), .A2(n717), .ZN(n515) );
  XNOR2_X1 U615 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n516) );
  XNOR2_X1 U616 ( .A(n517), .B(n516), .ZN(n729) );
  INV_X1 U617 ( .A(n518), .ZN(n519) );
  AND2_X1 U618 ( .A1(n701), .A2(n519), .ZN(n520) );
  INV_X1 U619 ( .A(n562), .ZN(n521) );
  NAND2_X1 U620 ( .A1(n561), .A2(n521), .ZN(n523) );
  INV_X1 U621 ( .A(KEYINPUT28), .ZN(n522) );
  INV_X1 U622 ( .A(n566), .ZN(n524) );
  INV_X1 U623 ( .A(KEYINPUT106), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n525), .B(KEYINPUT42), .ZN(n526) );
  XNOR2_X2 U625 ( .A(n527), .B(n526), .ZN(n672) );
  INV_X1 U626 ( .A(n672), .ZN(n528) );
  NAND2_X1 U627 ( .A1(n529), .A2(n528), .ZN(n532) );
  INV_X1 U628 ( .A(KEYINPUT84), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n530), .B(KEYINPUT46), .ZN(n531) );
  NAND2_X1 U630 ( .A1(n541), .A2(n535), .ZN(n755) );
  INV_X1 U631 ( .A(KEYINPUT73), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n718), .B(n536), .ZN(n538) );
  INV_X1 U633 ( .A(KEYINPUT47), .ZN(n537) );
  NAND2_X1 U634 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U635 ( .A1(n542), .A2(n378), .ZN(n546) );
  INV_X1 U636 ( .A(n543), .ZN(n576) );
  INV_X1 U637 ( .A(n544), .ZN(n613) );
  NOR2_X1 U638 ( .A1(n576), .A2(n613), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n677) );
  INV_X1 U640 ( .A(n718), .ZN(n554) );
  NAND2_X1 U641 ( .A1(n554), .A2(KEYINPUT47), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n677), .A2(n547), .ZN(n549) );
  INV_X1 U643 ( .A(KEYINPUT80), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U645 ( .A1(n677), .A2(KEYINPUT80), .ZN(n550) );
  NAND2_X1 U646 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U647 ( .A1(n554), .A2(KEYINPUT80), .ZN(n555) );
  NAND2_X1 U648 ( .A1(n555), .A2(n536), .ZN(n556) );
  NAND2_X1 U649 ( .A1(n557), .A2(KEYINPUT47), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U651 ( .A(n560), .B(KEYINPUT72), .ZN(n570) );
  XNOR2_X1 U652 ( .A(n705), .B(KEYINPUT6), .ZN(n616) );
  OR2_X1 U653 ( .A1(n574), .A2(n576), .ZN(n564) );
  INV_X1 U654 ( .A(KEYINPUT36), .ZN(n563) );
  XNOR2_X1 U655 ( .A(n564), .B(n563), .ZN(n568) );
  INV_X1 U656 ( .A(KEYINPUT1), .ZN(n565) );
  BUF_X1 U657 ( .A(n598), .Z(n567) );
  INV_X1 U658 ( .A(n567), .ZN(n699) );
  NAND2_X1 U659 ( .A1(n568), .A2(n699), .ZN(n757) );
  XNOR2_X1 U660 ( .A(n757), .B(KEYINPUT85), .ZN(n569) );
  INV_X1 U661 ( .A(KEYINPUT48), .ZN(n571) );
  INV_X1 U662 ( .A(n755), .ZN(n572) );
  NAND2_X1 U663 ( .A1(n573), .A2(n572), .ZN(n760) );
  OR2_X1 U664 ( .A1(n699), .A2(n574), .ZN(n575) );
  XNOR2_X1 U665 ( .A(n575), .B(KEYINPUT43), .ZN(n577) );
  NAND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n670) );
  AND2_X1 U667 ( .A1(n760), .A2(n670), .ZN(n578) );
  XNOR2_X1 U668 ( .A(KEYINPUT88), .B(G898), .ZN(n768) );
  NAND2_X1 U669 ( .A1(n768), .A2(G953), .ZN(n581) );
  AND2_X1 U670 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U671 ( .A1(n714), .A2(n586), .ZN(n587) );
  XOR2_X1 U672 ( .A(KEYINPUT100), .B(n587), .Z(n588) );
  XNOR2_X1 U673 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n589) );
  XNOR2_X1 U674 ( .A(n590), .B(n589), .ZN(n596) );
  OR2_X1 U675 ( .A1(n702), .A2(n567), .ZN(n591) );
  XNOR2_X1 U676 ( .A(n591), .B(KEYINPUT101), .ZN(n592) );
  AND2_X1 U677 ( .A1(n592), .A2(n616), .ZN(n593) );
  XOR2_X1 U678 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n594) );
  XNOR2_X1 U679 ( .A(n595), .B(n594), .ZN(n786) );
  AND2_X1 U680 ( .A1(n567), .A2(n596), .ZN(n619) );
  NOR2_X1 U681 ( .A1(n702), .A2(n705), .ZN(n597) );
  AND2_X1 U682 ( .A1(n619), .A2(n597), .ZN(n746) );
  INV_X1 U683 ( .A(n616), .ZN(n599) );
  INV_X1 U684 ( .A(KEYINPUT33), .ZN(n600) );
  XNOR2_X2 U685 ( .A(n601), .B(n600), .ZN(n712) );
  INV_X1 U686 ( .A(KEYINPUT70), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n603), .B(KEYINPUT34), .ZN(n604) );
  NOR2_X1 U688 ( .A1(n605), .A2(KEYINPUT44), .ZN(n608) );
  INV_X1 U689 ( .A(KEYINPUT44), .ZN(n606) );
  NOR2_X1 U690 ( .A1(n608), .A2(n607), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n678), .A2(KEYINPUT44), .ZN(n622) );
  INV_X1 U692 ( .A(n375), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n705), .A2(n610), .ZN(n708) );
  XNOR2_X1 U694 ( .A(n612), .B(KEYINPUT31), .ZN(n754) );
  NOR2_X1 U695 ( .A1(n613), .A2(n705), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n754), .A2(n743), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n615), .A2(n718), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n599), .A2(n617), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n673) );
  AND2_X1 U700 ( .A1(n620), .A2(n673), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(KEYINPUT86), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n629), .A2(KEYINPUT2), .ZN(n630) );
  INV_X1 U705 ( .A(n765), .ZN(n693) );
  INV_X1 U706 ( .A(n634), .ZN(n639) );
  NAND2_X1 U707 ( .A1(KEYINPUT2), .A2(n760), .ZN(n635) );
  XOR2_X1 U708 ( .A(KEYINPUT79), .B(n635), .Z(n637) );
  INV_X1 U709 ( .A(n670), .ZN(n636) );
  OR2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT83), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n374), .A2(G210), .ZN(n647) );
  XNOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n649) );
  INV_X1 U717 ( .A(G952), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n648), .A2(G953), .ZN(n690) );
  NAND2_X1 U719 ( .A1(n649), .A2(n690), .ZN(n651) );
  INV_X1 U720 ( .A(KEYINPUT56), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(G51) );
  NAND2_X1 U722 ( .A1(n374), .A2(G475), .ZN(n655) );
  XNOR2_X1 U723 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n656), .A2(n690), .ZN(n658) );
  INV_X1 U727 ( .A(KEYINPUT60), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(G60) );
  NAND2_X1 U729 ( .A1(n685), .A2(G478), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n661), .A2(n690), .ZN(n663) );
  INV_X1 U732 ( .A(KEYINPUT120), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G63) );
  NAND2_X1 U734 ( .A1(n685), .A2(G217), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n664), .B(KEYINPUT121), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n667), .A2(n690), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(G66) );
  XNOR2_X1 U739 ( .A(n670), .B(G140), .ZN(G42) );
  XNOR2_X1 U740 ( .A(G137), .B(KEYINPUT127), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(G39) );
  XNOR2_X1 U742 ( .A(n673), .B(G101), .ZN(G3) );
  XOR2_X1 U743 ( .A(G146), .B(KEYINPUT111), .Z(n676) );
  NOR2_X1 U744 ( .A1(n674), .A2(n751), .ZN(n675) );
  XOR2_X1 U745 ( .A(n676), .B(n675), .Z(G48) );
  XNOR2_X1 U746 ( .A(n677), .B(G143), .ZN(G45) );
  XOR2_X1 U747 ( .A(n376), .B(G122), .Z(G24) );
  NAND2_X1 U748 ( .A1(n374), .A2(G472), .ZN(n682) );
  XOR2_X1 U749 ( .A(KEYINPUT107), .B(KEYINPUT62), .Z(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n683), .A2(n690), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n684), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U754 ( .A1(n374), .A2(G469), .ZN(n689) );
  XOR2_X1 U755 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(n692) );
  INV_X1 U758 ( .A(n690), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(G54) );
  NOR2_X1 U760 ( .A1(n693), .A2(n780), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n694), .A2(KEYINPUT2), .ZN(n696) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n735) );
  NAND2_X1 U763 ( .A1(G952), .A2(n697), .ZN(n728) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U765 ( .A(KEYINPUT50), .B(n700), .Z(n707) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n703), .Z(n704) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U771 ( .A(n710), .B(KEYINPUT51), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n711), .A2(n729), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n719), .A2(n397), .ZN(n713) );
  XOR2_X1 U774 ( .A(KEYINPUT114), .B(n713), .Z(n716) );
  INV_X1 U775 ( .A(n714), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n722) );
  NAND2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n712), .A2(n723), .ZN(n724) );
  NOR2_X1 U781 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U782 ( .A(n726), .B(KEYINPUT52), .ZN(n727) );
  NOR2_X1 U783 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U784 ( .A1(n712), .A2(n729), .ZN(n730) );
  XOR2_X1 U785 ( .A(KEYINPUT115), .B(n730), .Z(n731) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U787 ( .A(KEYINPUT116), .B(n733), .Z(n734) );
  NOR2_X1 U788 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n736), .B(KEYINPUT117), .ZN(n737) );
  NOR2_X1 U790 ( .A1(n737), .A2(G953), .ZN(n739) );
  XNOR2_X1 U791 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n738) );
  XNOR2_X1 U792 ( .A(n739), .B(n738), .ZN(G75) );
  NOR2_X1 U793 ( .A1(n751), .A2(n743), .ZN(n740) );
  XOR2_X1 U794 ( .A(G104), .B(n740), .Z(G6) );
  XOR2_X1 U795 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n742) );
  XNOR2_X1 U796 ( .A(G107), .B(KEYINPUT108), .ZN(n741) );
  XNOR2_X1 U797 ( .A(n742), .B(n741), .ZN(n745) );
  NOR2_X1 U798 ( .A1(n755), .A2(n743), .ZN(n744) );
  XOR2_X1 U799 ( .A(n745), .B(n744), .Z(G9) );
  XNOR2_X1 U800 ( .A(G110), .B(n746), .ZN(n747) );
  XNOR2_X1 U801 ( .A(n747), .B(KEYINPUT109), .ZN(G12) );
  XOR2_X1 U802 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n749) );
  NOR2_X1 U803 ( .A1(n674), .A2(n755), .ZN(n748) );
  XOR2_X1 U804 ( .A(n749), .B(n748), .Z(n750) );
  XNOR2_X1 U805 ( .A(G128), .B(n750), .ZN(G30) );
  NOR2_X1 U806 ( .A1(n751), .A2(n754), .ZN(n752) );
  XOR2_X1 U807 ( .A(KEYINPUT112), .B(n752), .Z(n753) );
  XNOR2_X1 U808 ( .A(G113), .B(n753), .ZN(G15) );
  NOR2_X1 U809 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U810 ( .A(G116), .B(n756), .Z(G18) );
  XOR2_X1 U811 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n759) );
  XOR2_X1 U812 ( .A(G125), .B(n757), .Z(n758) );
  XNOR2_X1 U813 ( .A(n759), .B(n758), .ZN(G27) );
  XNOR2_X1 U814 ( .A(G134), .B(n760), .ZN(G36) );
  XOR2_X1 U815 ( .A(KEYINPUT125), .B(n761), .Z(n763) );
  NOR2_X1 U816 ( .A1(n768), .A2(n781), .ZN(n762) );
  NOR2_X1 U817 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U818 ( .A(KEYINPUT124), .B(n764), .ZN(n773) );
  NAND2_X1 U819 ( .A1(n765), .A2(n781), .ZN(n771) );
  XOR2_X1 U820 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n767) );
  NAND2_X1 U821 ( .A1(G224), .A2(G953), .ZN(n766) );
  XNOR2_X1 U822 ( .A(n767), .B(n766), .ZN(n769) );
  NAND2_X1 U823 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U824 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U825 ( .A(n773), .B(n772), .ZN(G69) );
  XNOR2_X1 U826 ( .A(n774), .B(n775), .ZN(n779) );
  XNOR2_X1 U827 ( .A(n779), .B(G227), .ZN(n776) );
  NAND2_X1 U828 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U829 ( .A1(G953), .A2(n777), .ZN(n778) );
  XNOR2_X1 U830 ( .A(n778), .B(KEYINPUT126), .ZN(n784) );
  XNOR2_X1 U831 ( .A(n780), .B(n779), .ZN(n782) );
  NAND2_X1 U832 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U833 ( .A1(n784), .A2(n783), .ZN(G72) );
  XOR2_X1 U834 ( .A(G131), .B(n785), .Z(G33) );
  XOR2_X1 U835 ( .A(G119), .B(n786), .Z(G21) );
endmodule

