//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0002(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n203));
  NAND2_X1  g0003(.A1(G116), .A2(G270), .ZN(new_n204));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  INV_X1    g0005(.A(G226), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n203), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n221), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n223), .A2(new_n230), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(G58), .A2(G68), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n219), .B1(new_n252), .B2(new_n205), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(G150), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n227), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n228), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n218), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n263), .B(new_n268), .C1(G50), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G222), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G223), .A2(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n282), .B(new_n285), .C1(G77), .C2(new_n278), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n218), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n289), .A2(G274), .A3(new_n284), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n287), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n286), .B(new_n291), .C1(new_n206), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g0095(.A(KEYINPUT72), .B(G200), .Z(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n272), .A2(new_n273), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n293), .A2(G179), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n293), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n270), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT75), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n206), .A2(new_n279), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n278), .B(new_n305), .C1(G232), .C2(new_n279), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n285), .ZN(new_n313));
  INV_X1    g0113(.A(new_n292), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G238), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n291), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n313), .A2(new_n318), .A3(new_n291), .A4(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(G190), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT12), .ZN(new_n321));
  INV_X1    g0121(.A(new_n269), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n269), .A2(KEYINPUT12), .A3(G68), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(new_n266), .B2(new_n323), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n275), .B1(new_n224), .B2(new_n226), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(G77), .B1(G50), .B2(new_n254), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n219), .B2(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n260), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT11), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n332), .A3(new_n260), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n326), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n320), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n317), .B2(new_n319), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n304), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n337), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n339), .A2(KEYINPUT75), .A3(new_n334), .A4(new_n320), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n317), .A2(new_n319), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(G169), .ZN(new_n344));
  AOI211_X1 g0144(.A(KEYINPUT14), .B(new_n301), .C1(new_n317), .C2(new_n319), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT76), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT76), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n317), .A2(new_n349), .A3(G179), .A4(new_n319), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n334), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT15), .B(G87), .Z(new_n354));
  NAND2_X1  g0154(.A1(new_n327), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT71), .ZN(new_n356));
  INV_X1    g0156(.A(G77), .ZN(new_n357));
  INV_X1    g0157(.A(new_n254), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n227), .A2(new_n357), .B1(new_n257), .B2(new_n358), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(KEYINPUT70), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n260), .B1(new_n357), .B2(new_n322), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n267), .A2(G77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G238), .A2(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n278), .B(new_n366), .C1(new_n212), .C2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n285), .C1(G107), .C2(new_n278), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n314), .A2(G244), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n291), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n296), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n370), .A2(new_n294), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n365), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n299), .A2(new_n303), .A3(new_n353), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n206), .A2(G1698), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n379), .B1(G223), .B2(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n284), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n291), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n292), .A2(new_n212), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n301), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n347), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n378), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(G179), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(KEYINPUT78), .C1(new_n387), .C2(new_n301), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT7), .B1(new_n278), .B2(G20), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n380), .A2(new_n381), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n227), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n394), .B(G68), .C1(KEYINPUT7), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(G58), .B(G68), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(new_n260), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n227), .A2(new_n395), .A3(KEYINPUT7), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n395), .B2(new_n219), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT77), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n227), .A2(new_n395), .A3(KEYINPUT77), .A4(KEYINPUT7), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n323), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n399), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n401), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n257), .A2(new_n269), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n267), .B2(new_n257), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n393), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n393), .A2(new_n414), .A3(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n387), .A2(new_n336), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT79), .B(G190), .Z(new_n421));
  NAND2_X1  g0221(.A1(new_n387), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n411), .A2(new_n420), .A3(new_n422), .A4(new_n413), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT17), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT73), .B1(new_n371), .B2(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G179), .B2(new_n370), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n371), .A2(KEYINPUT73), .A3(new_n347), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n365), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n419), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n377), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G250), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n276), .B2(new_n277), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n433));
  OAI211_X1 g0233(.A(G244), .B(new_n279), .C1(new_n380), .C2(new_n381), .ZN(new_n434));
  NOR2_X1   g0234(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT83), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT83), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n436), .A4(new_n433), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n285), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(G274), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n452), .A2(new_n284), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n449), .B1(new_n453), .B2(G257), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n444), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G200), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n269), .A2(G97), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n406), .A2(new_n407), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G107), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT6), .A2(G97), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n215), .A2(KEYINPUT80), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n460), .A2(new_n463), .A3(new_n465), .A4(new_n461), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n227), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n254), .A2(G77), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT81), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n227), .ZN(new_n473));
  INV_X1    g0273(.A(new_n468), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n463), .A2(new_n465), .B1(new_n460), .B2(new_n461), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n470), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n459), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n457), .B1(new_n479), .B2(new_n260), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n275), .A2(G1), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n322), .A2(new_n260), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G97), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n444), .A2(G190), .A3(new_n454), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n456), .A2(new_n480), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n472), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n215), .B1(new_n406), .B2(new_n407), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n260), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n457), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n483), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n455), .A2(new_n301), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n444), .A2(new_n347), .A3(new_n454), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  OR3_X1    g0294(.A1(new_n446), .A2(G1), .A3(G274), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n431), .B1(new_n446), .B2(G1), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n284), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OR2_X1    g0298(.A1(G238), .A2(G1698), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n278), .B(new_n499), .C1(G244), .C2(new_n279), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n285), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G190), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n285), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n497), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n296), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n309), .A2(KEYINPUT19), .A3(new_n310), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n227), .ZN(new_n511));
  NOR3_X1   g0311(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n256), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n227), .A2(new_n278), .A3(G68), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n354), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(new_n260), .B1(new_n322), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n482), .A2(G87), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n509), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(G169), .B1(new_n507), .B2(new_n497), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n482), .A2(new_n354), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n503), .A2(new_n347), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT84), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n503), .A2(new_n529), .A3(new_n347), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n506), .A2(new_n523), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n453), .A2(G264), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n431), .A2(new_n279), .ZN(new_n534));
  INV_X1    g0334(.A(G257), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n536), .C1(new_n380), .C2(new_n381), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n285), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n533), .A2(new_n540), .A3(new_n448), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT89), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n452), .A2(G264), .A3(new_n284), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n284), .B1(new_n537), .B2(new_n538), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(new_n449), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT89), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n547), .A3(new_n294), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(new_n336), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n227), .A2(new_n278), .A3(G87), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g0353(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n215), .A2(G20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(KEYINPUT23), .A2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n224), .A2(new_n226), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT22), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n227), .A2(new_n278), .A3(G87), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n553), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT24), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n553), .A2(new_n561), .A3(new_n567), .A4(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(new_n260), .B1(G107), .B2(new_n482), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n269), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n550), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n452), .A2(G270), .A3(new_n284), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT86), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n452), .A2(new_n576), .A3(G270), .A4(new_n284), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n449), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n279), .A2(G257), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n278), .B(new_n579), .C1(new_n216), .C2(new_n279), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n285), .C1(G303), .C2(new_n278), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n482), .A2(G116), .ZN(new_n583));
  INV_X1    g0383(.A(G116), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n322), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n275), .A2(G97), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n227), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n259), .A2(new_n228), .B1(G20), .B2(new_n584), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(KEYINPUT20), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT20), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n583), .B(new_n585), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n582), .A2(G169), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n582), .A2(G200), .ZN(new_n596));
  INV_X1    g0396(.A(new_n592), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n578), .A2(new_n421), .A3(new_n581), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n592), .A2(G179), .A3(new_n581), .A4(new_n578), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n582), .A2(KEYINPUT21), .A3(G169), .A4(new_n592), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n595), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n546), .A2(KEYINPUT89), .ZN(new_n603));
  NOR4_X1   g0403(.A1(new_n544), .A2(new_n545), .A3(new_n449), .A4(new_n542), .ZN(new_n604));
  OAI21_X1  g0404(.A(G169), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n546), .A2(G179), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n570), .A2(new_n572), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n573), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n430), .A2(new_n494), .A3(new_n532), .A4(new_n608), .ZN(G372));
  AOI21_X1  g0409(.A(KEYINPUT90), .B1(new_n526), .B2(new_n527), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n520), .A2(new_n322), .ZN(new_n611));
  INV_X1    g0411(.A(new_n518), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT19), .B1(new_n327), .B2(G97), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n512), .B1(new_n510), .B2(new_n227), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n611), .B(new_n525), .C1(new_n615), .C2(new_n264), .ZN(new_n616));
  INV_X1    g0416(.A(new_n524), .ZN(new_n617));
  AND4_X1   g0417(.A1(KEYINPUT90), .A2(new_n616), .A3(new_n617), .A4(new_n527), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(G169), .B1(new_n444), .B2(new_n454), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n444), .A2(new_n454), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n347), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n532), .A2(new_n622), .A3(new_n490), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n619), .B1(new_n623), .B2(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n616), .A2(new_n617), .A3(new_n527), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n509), .A2(new_n521), .A3(new_n504), .A4(new_n522), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n550), .A2(new_n570), .A3(new_n572), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n485), .B(new_n629), .C1(new_n607), .C2(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(KEYINPUT26), .B(new_n628), .C1(new_n631), .C2(new_n493), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n430), .B1(new_n625), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n391), .B1(new_n301), .B2(new_n387), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n414), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(new_n416), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n339), .A2(new_n334), .A3(new_n320), .ZN(new_n637));
  INV_X1    g0437(.A(new_n428), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n352), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT17), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n423), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n299), .B1(new_n270), .B2(new_n302), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n633), .A2(new_n643), .ZN(G369));
  OAI21_X1  g0444(.A(new_n629), .B1(new_n607), .B2(new_n630), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G13), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n473), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n218), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n655), .A2(new_n597), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n630), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n602), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n607), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n570), .A2(new_n572), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n664), .B(new_n629), .C1(new_n665), .C2(new_n655), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n630), .A2(new_n655), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n607), .A2(new_n654), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n658), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n231), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n513), .A2(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n229), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT92), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n655), .B1(new_n632), .B2(new_n625), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(KEYINPUT29), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n610), .B2(new_n618), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n626), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n526), .A2(KEYINPUT90), .A3(new_n527), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT94), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n532), .A2(new_n622), .A3(new_n690), .A4(new_n490), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT26), .B1(new_n493), .B2(new_n628), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n628), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n646), .A2(new_n493), .A3(new_n485), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n689), .A2(new_n691), .A3(new_n692), .A4(KEYINPUT95), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n682), .B1(new_n699), .B2(new_n655), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n681), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n608), .A2(new_n494), .A3(new_n532), .A4(new_n655), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n575), .A2(new_n577), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(G179), .A3(new_n448), .A4(new_n581), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n578), .A2(KEYINPUT93), .A3(G179), .A4(new_n581), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n533), .A2(new_n540), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n508), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n444), .A3(new_n454), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n703), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n707), .A2(new_n708), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n621), .A2(new_n714), .A3(KEYINPUT30), .A4(new_n711), .ZN(new_n715));
  AOI21_X1  g0515(.A(G179), .B1(new_n444), .B2(new_n454), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n508), .A3(new_n541), .A4(new_n582), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n702), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n718), .B2(new_n654), .ZN(new_n721));
  OAI21_X1  g0521(.A(G330), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n701), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n679), .B1(new_n723), .B2(G1), .ZN(G364));
  OR2_X1    g0524(.A1(new_n661), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n648), .A2(G45), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n674), .A2(G1), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT96), .Z(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n662), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n228), .B1(G20), .B2(new_n301), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n473), .A2(new_n294), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(G179), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G159), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n735), .A2(KEYINPUT32), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n372), .A2(G179), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(G20), .A3(G190), .ZN(new_n739));
  INV_X1    g0539(.A(G87), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n733), .A2(new_n372), .A3(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n278), .B1(new_n739), .B2(new_n740), .C1(new_n742), .C2(new_n215), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT97), .Z(new_n744));
  NAND3_X1  g0544(.A1(new_n347), .A2(new_n336), .A3(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n473), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G97), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT32), .B1(new_n735), .B2(new_n736), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n227), .A2(new_n347), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n748), .B1(new_n323), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n421), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n749), .A2(new_n336), .A3(new_n421), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n205), .B1(new_n758), .B2(new_n211), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n744), .A2(new_n747), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n749), .A2(new_n294), .A3(new_n336), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n737), .B(new_n761), .C1(G77), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n734), .A2(G329), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n752), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n742), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G322), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n758), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n768), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n739), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G303), .B1(G294), .B2(new_n746), .ZN(new_n775));
  AND3_X1   g0575(.A1(new_n773), .A2(new_n395), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n776), .B1(new_n777), .B2(new_n762), .C1(new_n778), .C2(new_n756), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n732), .B1(new_n765), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n231), .A2(G355), .A3(new_n278), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n672), .A2(new_n278), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G45), .B2(new_n229), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n247), .A2(new_n446), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n781), .B1(G116), .B2(new_n231), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n731), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n728), .B(new_n790), .C1(new_n661), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n730), .B1(new_n780), .B2(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n731), .A2(new_n786), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n729), .B1(new_n357), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n365), .A2(new_n654), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n428), .B1(new_n375), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n638), .A2(new_n655), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n751), .A2(G150), .B1(new_n757), .B2(G143), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n756), .C1(new_n736), .C2(new_n762), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n741), .A2(G68), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n395), .B1(new_n746), .B2(G58), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n205), .B2(new_n739), .C1(new_n808), .C2(new_n735), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n774), .A2(G107), .B1(G116), .B2(new_n763), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n777), .B2(new_n735), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n758), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n752), .A2(new_n769), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n741), .A2(G87), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n755), .A2(G303), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n815), .A2(new_n747), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n809), .B1(new_n278), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT99), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n795), .B1(new_n787), .B2(new_n800), .C1(new_n820), .C2(new_n732), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n680), .A2(new_n799), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n655), .B(new_n800), .C1(new_n632), .C2(new_n625), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n722), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n729), .B1(new_n824), .B2(new_n722), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT101), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  NOR2_X1   g0630(.A1(new_n474), .A2(new_n475), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT102), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT35), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n228), .B(new_n227), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(G116), .C1(new_n833), .C2(new_n832), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  OAI21_X1  g0636(.A(G77), .B1(new_n211), .B2(new_n323), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n229), .B1(G50), .B2(new_n323), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(G1), .A3(new_n647), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT103), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n655), .A2(new_n334), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n341), .B2(new_n352), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n346), .A2(new_n351), .ZN(new_n844));
  INV_X1    g0644(.A(new_n334), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n842), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n847), .A2(new_n637), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n400), .A2(new_n260), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT16), .B1(new_n397), .B2(new_n399), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n413), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n652), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n419), .B2(new_n424), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n634), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n423), .A2(new_n858), .A3(new_n856), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n414), .A2(new_n855), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n415), .A2(new_n861), .A3(new_n862), .A4(new_n423), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n851), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n856), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n393), .A2(new_n414), .A3(KEYINPUT18), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT18), .B1(new_n393), .B2(new_n414), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n866), .B1(new_n869), .B2(new_n641), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n860), .A2(new_n863), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n872));
  AOI221_X4 g0672(.A(new_n850), .B1(new_n865), .B2(new_n872), .C1(new_n823), .C2(new_n798), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n636), .A2(new_n855), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT104), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n865), .A2(new_n872), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n861), .B1(new_n636), .B2(new_n424), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n635), .A2(new_n861), .A3(new_n423), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n863), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n851), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n872), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n846), .A2(new_n654), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n878), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n850), .ZN(new_n889));
  INV_X1    g0689(.A(new_n485), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n493), .B1(new_n645), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n690), .A3(new_n696), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n654), .B(new_n799), .C1(new_n892), .C2(new_n624), .ZN(new_n893));
  INV_X1    g0693(.A(new_n798), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n876), .B(new_n889), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT104), .ZN(new_n896));
  INV_X1    g0696(.A(new_n874), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n875), .A2(new_n888), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n430), .B1(new_n700), .B2(new_n681), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n643), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n899), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT105), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n718), .A2(new_n904), .A3(new_n654), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT31), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n904), .B1(new_n718), .B2(new_n654), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n719), .B(new_n702), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n799), .B1(new_n843), .B2(new_n849), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n903), .B1(new_n877), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n910), .A4(new_n909), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n912), .A2(new_n913), .A3(new_n909), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(G330), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n430), .A2(G330), .A3(new_n909), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n914), .A2(new_n430), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n902), .B(new_n917), .Z(new_n918));
  NOR2_X1   g0718(.A1(new_n648), .A2(new_n218), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n841), .B1(new_n918), .B2(new_n919), .ZN(G367));
  AOI21_X1  g0720(.A(new_n655), .B1(new_n521), .B2(new_n522), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n921), .A2(new_n628), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n619), .A2(new_n921), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n729), .B1(new_n925), .B2(new_n788), .ZN(new_n926));
  INV_X1    g0726(.A(new_n782), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n789), .B1(new_n231), .B2(new_n520), .C1(new_n243), .C2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(G97), .A2(new_n741), .B1(new_n763), .B2(G283), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n739), .A2(new_n584), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n929), .B1(new_n777), .B2(new_n756), .C1(new_n930), .C2(KEYINPUT46), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(KEYINPUT46), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n812), .B2(new_n752), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n278), .B(new_n933), .C1(G317), .C2(new_n734), .ZN(new_n934));
  INV_X1    g0734(.A(new_n746), .ZN(new_n935));
  INV_X1    g0735(.A(G303), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n934), .B1(new_n215), .B2(new_n935), .C1(new_n936), .C2(new_n758), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n323), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n741), .A2(G77), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n939), .B1(new_n739), .B2(new_n211), .C1(new_n752), .C2(new_n736), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G143), .B2(new_n755), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n278), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n938), .B(new_n942), .C1(G137), .C2(new_n734), .ZN(new_n943));
  INV_X1    g0743(.A(G150), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(new_n205), .B2(new_n762), .C1(new_n944), .C2(new_n758), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n937), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  OAI211_X1 g0747(.A(new_n926), .B(new_n928), .C1(new_n947), .C2(new_n732), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n726), .A2(G1), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n490), .A2(new_n654), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n494), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n622), .A2(new_n490), .A3(new_n654), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n658), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT44), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n658), .A2(new_n953), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT45), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n670), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n663), .A2(new_n669), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n664), .A2(new_n629), .A3(new_n630), .A4(new_n655), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n670), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n723), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n723), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n673), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n949), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n670), .B1(new_n951), .B2(new_n952), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n925), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(KEYINPUT109), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT108), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n493), .B1(new_n951), .B2(new_n664), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT107), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n655), .ZN(new_n980));
  INV_X1    g0780(.A(new_n494), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n962), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n977), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n973), .A2(KEYINPUT109), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n975), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n984), .A2(KEYINPUT109), .A3(new_n973), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n971), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n970), .A3(new_n987), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n948), .B1(new_n969), .B2(new_n993), .ZN(G387));
  NOR2_X1   g0794(.A1(new_n723), .A2(new_n964), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT114), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n965), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n673), .C1(new_n996), .C2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n675), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n257), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(G68), .A2(G77), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n257), .B2(G50), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1001), .A2(new_n446), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n782), .B(new_n1004), .C1(new_n239), .C2(new_n446), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n999), .A2(new_n231), .A3(new_n278), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G107), .C2(new_n231), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT110), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n789), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n739), .A2(new_n357), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n752), .A2(new_n257), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n758), .A2(new_n205), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n935), .A2(new_n520), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n323), .B2(new_n762), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1010), .B(new_n1015), .C1(G150), .C2(new_n734), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n736), .B2(new_n756), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n395), .B(new_n1017), .C1(G97), .C2(new_n741), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n751), .A2(G311), .B1(new_n757), .B2(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n936), .B2(new_n762), .C1(new_n771), .C2(new_n756), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n739), .A2(new_n812), .B1(new_n769), .B2(new_n935), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT111), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  OAI221_X1 g0827(.A(new_n395), .B1(new_n735), .B2(new_n778), .C1(new_n742), .C2(new_n584), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(KEYINPUT112), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(KEYINPUT112), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1018), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n728), .B(new_n1009), .C1(new_n1032), .C2(new_n732), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT113), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n666), .A2(new_n668), .A3(new_n788), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n949), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n998), .B(new_n1036), .C1(new_n1037), .C2(new_n963), .ZN(G393));
  OR2_X1    g0838(.A1(new_n959), .A2(new_n670), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(new_n960), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n673), .B(new_n966), .C1(new_n1040), .C2(new_n965), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n949), .A3(new_n960), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n789), .B1(new_n927), .B2(new_n250), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G97), .B2(new_n672), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n755), .A2(G150), .B1(new_n757), .B2(G159), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n278), .B1(new_n762), .B2(new_n257), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n816), .B1(new_n752), .B2(new_n205), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n774), .A2(G68), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n734), .A2(G143), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1045), .A2(KEYINPUT51), .B1(G77), .B2(new_n746), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n755), .A2(G317), .B1(new_n757), .B2(G311), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n278), .B(new_n1055), .C1(G322), .C2(new_n734), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n751), .A2(G303), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n763), .A2(G294), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n741), .A2(G107), .B1(G116), .B2(new_n746), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n739), .A2(new_n769), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1053), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n729), .B(new_n1044), .C1(new_n1062), .C2(new_n731), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n791), .B2(new_n953), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1042), .A2(KEYINPUT115), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(KEYINPUT115), .B1(new_n1042), .B2(new_n1064), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1041), .B1(new_n1065), .B2(new_n1066), .ZN(G390));
  NAND3_X1  g0867(.A1(new_n699), .A2(new_n655), .A3(new_n797), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n798), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT116), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(KEYINPUT116), .A3(new_n798), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n889), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n887), .B1(new_n883), .B2(new_n872), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n878), .A2(new_n886), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n850), .B1(new_n823), .B2(new_n798), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(new_n887), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1073), .A2(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n722), .A2(new_n799), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n889), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n909), .A2(new_n910), .A3(G330), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT117), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT117), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n909), .A2(new_n910), .A3(new_n1085), .A4(G330), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1082), .B1(new_n1087), .B2(new_n1078), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1079), .A2(new_n889), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1087), .A2(new_n1090), .B1(new_n894), .B2(new_n893), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n907), .A2(new_n908), .ZN(new_n1092));
  OAI211_X1 g0892(.A(G330), .B(new_n800), .C1(new_n1092), .C2(new_n720), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n850), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(KEYINPUT118), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT118), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n1096), .A3(new_n850), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1068), .A2(KEYINPUT116), .A3(new_n798), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT116), .B1(new_n1068), .B2(new_n798), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1095), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1091), .B1(new_n1100), .B2(new_n1081), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT119), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n900), .A2(new_n916), .A3(new_n643), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1102), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT120), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT119), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT120), .B1(new_n1111), .B2(new_n1105), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1089), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1088), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n673), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1089), .A2(new_n1037), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n755), .A2(G128), .B1(new_n757), .B2(G132), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT121), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G50), .B2(new_n741), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n746), .A2(G159), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT54), .B(G143), .Z(new_n1121));
  NAND2_X1  g0921(.A1(new_n763), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n752), .B2(new_n802), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n395), .B(new_n1123), .C1(G125), .C2(new_n734), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n739), .A2(new_n944), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT53), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1119), .A2(new_n1120), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n805), .B1(new_n735), .B2(new_n812), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT122), .Z(new_n1129));
  OAI22_X1  g0929(.A1(new_n756), .A2(new_n769), .B1(new_n758), .B2(new_n584), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n395), .B1(new_n935), .B2(new_n357), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n739), .A2(new_n740), .B1(new_n516), .B2(new_n762), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1129), .B(new_n1133), .C1(new_n215), .C2(new_n752), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n732), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n729), .B(new_n1135), .C1(new_n257), .C2(new_n794), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1075), .B2(new_n786), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1116), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1115), .A2(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1111), .A2(new_n1105), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1103), .B1(new_n1142), .B2(new_n1088), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n299), .A2(new_n303), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1145));
  XOR2_X1   g0945(.A(new_n1144), .B(new_n1145), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n270), .A2(new_n855), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(KEYINPUT104), .B(new_n874), .C1(new_n1076), .C2(new_n876), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n915), .B1(new_n1152), .B2(new_n888), .ZN(new_n1153));
  AND4_X1   g0953(.A1(new_n915), .A2(new_n875), .A3(new_n888), .A4(new_n898), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n915), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n899), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1152), .A2(new_n915), .A3(new_n888), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1148), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1141), .B1(new_n1143), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1114), .A2(new_n1104), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1160), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(KEYINPUT57), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1164), .A3(new_n673), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1155), .A2(new_n949), .A3(new_n1159), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n794), .A2(new_n205), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n742), .A2(new_n211), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n516), .A2(new_n752), .B1(new_n756), .B2(new_n584), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n354), .C2(new_n763), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n395), .B1(new_n735), .B2(new_n769), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1171), .A2(new_n1010), .A3(G41), .A4(new_n938), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n215), .C2(new_n758), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT58), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n205), .B1(new_n380), .B2(G41), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n774), .A2(new_n1121), .B1(G128), .B2(new_n757), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n746), .A2(G150), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G125), .A2(new_n755), .B1(new_n763), .B2(G137), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G132), .B2(new_n751), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT59), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G33), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G41), .B1(new_n734), .B2(G124), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n736), .C2(new_n742), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1174), .B(new_n1175), .C1(new_n1182), .C2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT123), .Z(new_n1187));
  AOI21_X1  g0987(.A(new_n729), .B1(new_n1187), .B2(new_n731), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1167), .B(new_n1188), .C1(new_n1148), .C2(new_n787), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1166), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(G375));
  OAI21_X1  g0992(.A(new_n1108), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1111), .A2(KEYINPUT120), .A3(new_n1105), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n968), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1101), .A2(new_n949), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G294), .A2(new_n755), .B1(new_n763), .B2(G107), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n516), .B2(new_n739), .C1(new_n584), .C2(new_n752), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G283), .B2(new_n757), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n278), .B(new_n1013), .C1(new_n734), .C2(G303), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n939), .A3(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT124), .Z(new_n1205));
  AOI22_X1  g1005(.A1(new_n751), .A2(new_n1121), .B1(new_n763), .B2(G150), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1206), .B(new_n278), .C1(new_n736), .C2(new_n739), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n935), .A2(new_n205), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n734), .A2(G128), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1207), .A2(new_n1168), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n808), .B2(new_n756), .C1(new_n802), .C2(new_n758), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n732), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n729), .B(new_n1212), .C1(new_n323), .C2(new_n794), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n787), .B2(new_n889), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1199), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1198), .A2(new_n1216), .ZN(G381));
  AOI21_X1  g1017(.A(new_n1160), .B1(new_n1114), .B2(new_n1104), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n674), .B1(new_n1218), .B2(KEYINPUT57), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1190), .B1(new_n1219), .B2(new_n1161), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1139), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1114), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1195), .B2(new_n1089), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1221), .B1(new_n1223), .B2(new_n673), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G384), .A3(G381), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G390), .A2(G387), .ZN(new_n1227));
  OR2_X1    g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1229), .ZN(G407));
  OAI211_X1 g1030(.A(G407), .B(G213), .C1(G343), .C2(new_n1225), .ZN(G409));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1218), .A2(new_n968), .B1(new_n1190), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1191), .A2(KEYINPUT125), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1233), .A2(new_n1115), .A3(new_n1139), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n653), .A2(G213), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G375), .A2(G378), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1101), .A2(new_n1104), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n1105), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n674), .B(new_n1240), .C1(new_n1241), .C2(new_n1197), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n829), .B1(new_n1242), .B2(new_n1215), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1197), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1240), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n673), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(G384), .A3(new_n1216), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n653), .A2(KEYINPUT126), .A3(G213), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1243), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1250), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1243), .A2(new_n1247), .A3(new_n1252), .A4(new_n1248), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1237), .A2(new_n1238), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1235), .B(new_n1236), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT63), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1256), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1238), .A2(new_n1259), .A3(new_n1236), .A4(new_n1235), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1228), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1227), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G390), .A2(G387), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(G390), .A2(G387), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1228), .B(new_n1263), .C1(new_n1268), .C2(new_n1227), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT127), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1258), .A2(new_n1262), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1255), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT62), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1270), .B1(new_n1260), .B2(KEYINPUT62), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1274), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1280), .ZN(G405));
  NAND2_X1  g1081(.A1(new_n1238), .A2(new_n1225), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1269), .A3(new_n1267), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1274), .A2(new_n1225), .A3(new_n1238), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1259), .ZN(G402));
endmodule


