//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n208), .A3(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT88), .ZN(new_n212));
  AND2_X1   g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G43gat), .A2(G50gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT15), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT14), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT14), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G29gat), .B2(G36gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n212), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n231), .A2(KEYINPUT88), .A3(new_n215), .A4(new_n221), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  INV_X1    g033(.A(new_n215), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT87), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n228), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT87), .B1(new_n225), .B2(new_n227), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n233), .A2(new_n234), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n234), .B1(new_n233), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n211), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT90), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n210), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n233), .A2(new_n239), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n207), .A2(KEYINPUT90), .A3(new_n209), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT89), .B(new_n211), .C1(new_n240), .C2(new_n241), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n244), .A2(new_n245), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(G229gat), .B2(G233gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n244), .A2(new_n250), .A3(new_n251), .A4(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n233), .A2(new_n239), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n207), .A2(KEYINPUT90), .A3(new_n209), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT90), .B1(new_n207), .B2(new_n209), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n250), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n245), .B(KEYINPUT13), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n254), .A2(new_n256), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G169gat), .B(G197gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT12), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n252), .A2(new_n253), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n261), .B2(new_n262), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n256), .A2(new_n274), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT91), .B1(new_n278), .B2(new_n254), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n272), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G148gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT79), .B(G141gat), .Z(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  OR2_X1    g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(KEYINPUT2), .ZN(new_n288));
  XNOR2_X1  g087(.A(G141gat), .B(G148gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(KEYINPUT2), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n285), .A2(new_n288), .B1(new_n290), .B2(KEYINPUT78), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n287), .A2(new_n286), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n292), .B(new_n293), .C1(KEYINPUT2), .C2(new_n289), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT71), .B(G134gat), .C1(new_n295), .C2(KEYINPUT1), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G127gat), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n296), .B2(new_n303), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n291), .B(new_n294), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n285), .A2(new_n288), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n290), .A2(KEYINPUT78), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n294), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n305), .B2(new_n306), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n301), .A2(new_n316), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n295), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n318));
  OAI21_X1  g117(.A(G127gat), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT80), .A4(new_n294), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n313), .A2(new_n315), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n308), .B1(new_n323), .B2(KEYINPUT4), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n305), .A2(new_n306), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n291), .A2(new_n327), .A3(new_n294), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(KEYINPUT84), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n326), .A2(new_n311), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n307), .A3(new_n331), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n335), .A2(KEYINPUT39), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT39), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT84), .B1(new_n330), .B2(new_n332), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n334), .B(new_n331), .C1(new_n324), .C2(new_n329), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT85), .ZN(new_n344));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT0), .ZN(new_n346));
  XNOR2_X1  g145(.A(G57gat), .B(G85gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n344), .B1(new_n343), .B2(new_n348), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n339), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT40), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n307), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n332), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n357), .B2(KEYINPUT81), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n359), .A3(new_n332), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n323), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n307), .A2(new_n361), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n329), .A2(new_n363), .A3(new_n331), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n358), .B(new_n360), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n324), .A2(new_n355), .A3(new_n331), .A4(new_n329), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n348), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(G197gat), .A2(G204gat), .ZN(new_n368));
  AND2_X1   g167(.A1(G197gat), .A2(G204gat), .ZN(new_n369));
  AND2_X1   g168(.A1(G211gat), .A2(G218gat), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n368), .A2(new_n369), .B1(new_n370), .B2(KEYINPUT22), .ZN(new_n371));
  XOR2_X1   g170(.A(G211gat), .B(G218gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G226gat), .ZN(new_n374));
  INV_X1    g173(.A(G233gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(KEYINPUT24), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(KEYINPUT67), .ZN(new_n383));
  OAI221_X1 g182(.A(new_n378), .B1(G183gat), .B2(G190gat), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n385));
  INV_X1    g184(.A(G169gat), .ZN(new_n386));
  INV_X1    g185(.A(G176gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(KEYINPUT65), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  NOR2_X1   g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(KEYINPUT23), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n385), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT66), .B1(new_n395), .B2(new_n396), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n384), .B(new_n394), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n402));
  INV_X1    g201(.A(new_n397), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(new_n393), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n406));
  OAI221_X1 g205(.A(new_n378), .B1(G183gat), .B2(G190gat), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n403), .B(new_n404), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n401), .A2(new_n402), .B1(new_n385), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n397), .B(new_n398), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n411), .A2(KEYINPUT68), .A3(new_n384), .A4(new_n394), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT27), .B(G183gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT69), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G190gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT28), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n413), .A2(new_n416), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n418), .A2(KEYINPUT28), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n388), .A2(KEYINPUT26), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT70), .ZN(new_n422));
  INV_X1    g221(.A(new_n396), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(KEYINPUT26), .B2(new_n388), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n422), .A2(new_n424), .B1(G183gat), .B2(G190gat), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n410), .A2(new_n412), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n377), .B1(new_n426), .B2(KEYINPUT29), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n426), .A2(new_n428), .A3(new_n377), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n401), .A2(new_n402), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n385), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n420), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT75), .B1(new_n434), .B2(new_n376), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n373), .B(new_n427), .C1(new_n429), .C2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n373), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n376), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n426), .A2(new_n377), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G64gat), .B(G92gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n436), .A2(new_n441), .ZN(new_n448));
  INV_X1    g247(.A(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n445), .A2(KEYINPUT76), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT76), .B1(new_n445), .B2(new_n452), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n367), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n343), .A2(new_n348), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT85), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n349), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(KEYINPUT40), .A3(new_n339), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n354), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n436), .A2(new_n441), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n444), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT38), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n437), .B(new_n427), .C1(new_n429), .C2(new_n435), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n373), .B1(new_n439), .B2(new_n440), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT37), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n357), .A2(KEYINPUT81), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT5), .A3(new_n360), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n362), .A2(new_n364), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n348), .B(new_n366), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n367), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n366), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  INV_X1    g276(.A(new_n348), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n474), .A3(new_n473), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n469), .A2(new_n476), .A3(new_n480), .A4(new_n445), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n448), .A2(KEYINPUT37), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n465), .B1(new_n464), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n373), .B1(new_n328), .B2(new_n438), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n313), .A2(new_n322), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n371), .A2(KEYINPUT82), .A3(new_n372), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n438), .B(new_n490), .C1(new_n373), .C2(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n327), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n311), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT3), .B1(new_n373), .B2(new_n438), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n486), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(new_n487), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G78gat), .B(G106gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT31), .B(G50gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n502), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n494), .B2(new_n498), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n506));
  INV_X1    g305(.A(G22gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n505), .B2(new_n506), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n488), .A2(new_n493), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n485), .ZN(new_n513));
  INV_X1    g312(.A(new_n498), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(G22gat), .B1(new_n515), .B2(KEYINPUT83), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n516), .A2(new_n502), .A3(new_n499), .A4(new_n508), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n461), .A2(new_n484), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G227gat), .A2(G233gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n315), .A2(new_n321), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n434), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n315), .A2(new_n321), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n426), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT32), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G15gat), .B(G43gat), .Z(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n434), .A2(new_n523), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n426), .A2(new_n525), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n521), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT34), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n521), .B1(new_n535), .B2(new_n536), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n540), .B2(KEYINPUT33), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT32), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n534), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT73), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n534), .A2(new_n544), .A3(new_n547), .A4(new_n539), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n537), .B(KEYINPUT34), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n541), .A2(new_n543), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n536), .ZN(new_n551));
  AOI221_X4 g350(.A(new_n542), .B1(KEYINPUT33), .B2(new_n533), .C1(new_n551), .C2(new_n522), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n544), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n549), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n546), .B(new_n548), .C1(new_n554), .C2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(KEYINPUT36), .A3(new_n545), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n480), .A2(new_n476), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n454), .A2(new_n562), .A3(new_n455), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n560), .A2(new_n561), .B1(new_n518), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n520), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n475), .B(new_n479), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n462), .A2(new_n567), .A3(KEYINPUT30), .A4(new_n444), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n568), .A2(new_n455), .A3(new_n447), .A4(new_n450), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n555), .A3(new_n549), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n511), .A2(new_n517), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n546), .A2(new_n548), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n573), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n511), .A2(new_n517), .A3(new_n553), .A4(new_n545), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT35), .B1(new_n563), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n281), .B1(new_n565), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT96), .ZN(new_n584));
  XOR2_X1   g383(.A(G134gat), .B(G162gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n591), .A2(new_n592), .B1(KEYINPUT8), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT97), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n595), .A2(new_n597), .A3(G85gat), .A4(G92gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G92gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n594), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n594), .A2(new_n598), .A3(new_n606), .A4(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n589), .B1(new_n257), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT99), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n240), .B2(new_n241), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n587), .B(new_n588), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n616), .A2(new_n587), .A3(new_n618), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G57gat), .B(G64gat), .Z(new_n623));
  INV_X1    g422(.A(KEYINPUT9), .ZN(new_n624));
  INV_X1    g423(.A(G71gat), .ZN(new_n625));
  INV_X1    g424(.A(G78gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G71gat), .B(G78gat), .ZN(new_n629));
  OR2_X1    g428(.A1(G57gat), .A2(G64gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n631));
  NAND2_X1  g430(.A1(G57gat), .A2(G64gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n627), .A3(new_n623), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n634), .A2(new_n636), .A3(KEYINPUT95), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT21), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n258), .B2(new_n259), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT93), .B(KEYINPUT94), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n647));
  AND2_X1   g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G183gat), .B(G211gat), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n655), .B1(new_n652), .B2(new_n653), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n646), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n645), .A3(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n610), .A2(new_n637), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n608), .A2(new_n636), .A3(new_n634), .A4(new_n609), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT10), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n639), .B2(new_n640), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n669), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(new_n668), .A3(new_n671), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G120gat), .B(G148gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT101), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n622), .A2(new_n667), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n582), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n562), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(G1gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1324gat));
  XNOR2_X1  g489(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n208), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n582), .A2(new_n569), .A3(new_n686), .A4(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n582), .A2(new_n569), .A3(new_n686), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G8gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n693), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(KEYINPUT42), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT104), .ZN(G1325gat));
  AOI21_X1  g499(.A(KEYINPUT36), .B1(new_n577), .B2(new_n573), .ZN(new_n701));
  INV_X1    g500(.A(new_n561), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n687), .B2(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n558), .A2(G15gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n687), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n687), .A2(new_n519), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n667), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n685), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n622), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT105), .Z(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(new_n582), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n223), .A3(new_n566), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n558), .A2(new_n563), .A3(new_n575), .ZN(new_n719));
  INV_X1    g518(.A(new_n579), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n574), .B1(new_n570), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n578), .A2(new_n723), .A3(new_n580), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n722), .A2(new_n724), .B1(new_n520), .B2(new_n564), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n718), .B1(new_n725), .B2(new_n622), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n565), .A2(new_n581), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(KEYINPUT44), .A3(new_n621), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n276), .B1(new_n273), .B2(new_n275), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n278), .A2(KEYINPUT91), .A3(new_n254), .ZN(new_n730));
  AOI221_X4 g529(.A(KEYINPUT106), .B1(new_n264), .B2(new_n271), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n272), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n712), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n726), .A2(new_n728), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n562), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n717), .A2(new_n739), .ZN(G1328gat));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  AOI21_X1  g540(.A(G36gat), .B1(new_n741), .B2(KEYINPUT46), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n715), .A2(new_n569), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n569), .ZN(new_n746));
  OAI21_X1  g545(.A(G36gat), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1329gat));
  OAI21_X1  g547(.A(G43gat), .B1(new_n738), .B2(new_n704), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT47), .B1(new_n749), .B2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g549(.A(new_n558), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n715), .A2(new_n216), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n749), .B(new_n752), .C1(KEYINPUT109), .C2(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1330gat));
  OAI21_X1  g555(.A(G50gat), .B1(new_n738), .B2(new_n519), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n715), .A2(new_n217), .A3(new_n518), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1331gat));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n736), .A2(new_n667), .A3(new_n622), .A4(new_n684), .ZN(new_n763));
  OR3_X1    g562(.A1(new_n725), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n725), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n566), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n569), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT49), .B(G64gat), .Z(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n766), .B2(new_n704), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n764), .A2(new_n765), .A3(new_n625), .A4(new_n751), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(KEYINPUT50), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n766), .A2(new_n519), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n626), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n735), .A2(new_n667), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n684), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n726), .A2(new_n728), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n562), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n578), .A2(new_n723), .A3(new_n580), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n723), .B1(new_n578), .B2(new_n580), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n519), .B1(new_n481), .B2(new_n483), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT40), .B1(new_n459), .B2(new_n339), .ZN(new_n791));
  INV_X1    g590(.A(new_n339), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n353), .B(new_n792), .C1(new_n458), .C2(new_n349), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n794), .B2(new_n456), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n701), .A2(new_n702), .B1(new_n519), .B2(new_n570), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n788), .A2(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n621), .A3(new_n783), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n797), .A2(new_n800), .A3(new_n621), .A4(new_n783), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n684), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n566), .A2(new_n603), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n787), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NAND4_X1  g603(.A1(new_n726), .A2(new_n569), .A3(new_n728), .A4(new_n785), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n600), .A2(new_n602), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n746), .A2(G92gat), .A3(new_n685), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n810), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n621), .A3(new_n783), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n807), .B1(new_n814), .B2(KEYINPUT113), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n801), .A3(new_n808), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n807), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1337gat));
  OAI21_X1  g620(.A(G99gat), .B1(new_n786), .B2(new_n704), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n558), .A2(G99gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n799), .A2(new_n684), .A3(new_n801), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT114), .ZN(G1338gat));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n813), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n519), .A2(G106gat), .A3(new_n685), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n726), .A2(new_n518), .A3(new_n728), .A4(new_n785), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT53), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n799), .A2(new_n801), .A3(new_n828), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT115), .B1(new_n836), .B2(new_n831), .ZN(new_n837));
  AND4_X1   g636(.A1(KEYINPUT115), .A2(new_n831), .A3(new_n835), .A4(new_n834), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(G1339gat));
  AND2_X1   g638(.A1(new_n251), .A2(new_n250), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n245), .B1(new_n840), .B2(new_n244), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n841), .A2(KEYINPUT119), .B1(new_n261), .B2(new_n262), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n269), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n733), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n672), .A2(new_n674), .A3(new_n669), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n675), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n669), .C1(new_n672), .C2(new_n674), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(KEYINPUT117), .A3(new_n681), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n851), .B2(new_n681), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n851), .A2(new_n681), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n851), .A2(KEYINPUT117), .A3(new_n681), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n849), .ZN(new_n863));
  AND4_X1   g662(.A1(new_n682), .A2(new_n856), .A3(new_n857), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n864), .A3(new_n621), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n845), .A2(new_n733), .A3(new_n684), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n735), .B2(new_n864), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT120), .B(new_n865), .C1(new_n867), .C2(new_n621), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n280), .A2(KEYINPUT106), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n733), .A2(new_n732), .A3(new_n272), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n864), .ZN(new_n872));
  INV_X1    g671(.A(new_n866), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n621), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n865), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n876), .A3(new_n711), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n686), .A2(KEYINPUT116), .A3(new_n736), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT116), .B1(new_n686), .B2(new_n736), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n518), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n569), .A2(new_n562), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n751), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n299), .A3(new_n281), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n877), .A2(new_n880), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n882), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n720), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n735), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(new_n299), .ZN(G1340gat));
  NOR3_X1   g688(.A1(new_n883), .A2(new_n297), .A3(new_n685), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n684), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n297), .ZN(G1341gat));
  XOR2_X1   g691(.A(KEYINPUT71), .B(G127gat), .Z(new_n893));
  NOR3_X1   g692(.A1(new_n883), .A2(new_n711), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n887), .A2(new_n667), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n893), .ZN(G1342gat));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n622), .A2(G134gat), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n886), .A2(new_n897), .A3(new_n720), .A4(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT121), .ZN(new_n900));
  OAI21_X1  g699(.A(G134gat), .B1(new_n883), .B2(new_n622), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n887), .A2(new_n898), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n900), .B(new_n901), .C1(new_n897), .C2(new_n902), .ZN(G1343gat));
  NOR2_X1   g702(.A1(new_n703), .A2(new_n519), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n281), .A2(G141gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n857), .B(KEYINPUT122), .Z(new_n909));
  AND3_X1   g708(.A1(new_n856), .A2(new_n682), .A3(new_n863), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n280), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n621), .B1(new_n911), .B2(new_n873), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n711), .B1(new_n912), .B2(new_n875), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n880), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n518), .A2(KEYINPUT57), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n519), .B1(new_n877), .B2(new_n880), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(KEYINPUT57), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n703), .A2(new_n562), .A3(new_n569), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n280), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n919), .A2(KEYINPUT123), .A3(new_n280), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n284), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n908), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n885), .B2(new_n518), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n915), .B1(new_n880), .B2(new_n913), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n735), .B(new_n920), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n284), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n906), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(new_n932), .ZN(G1344gat));
  NAND2_X1  g732(.A1(new_n919), .A2(new_n920), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n934), .A2(KEYINPUT59), .A3(new_n685), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n886), .A2(new_n904), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT59), .B1(new_n936), .B2(new_n685), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n282), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n915), .B1(new_n877), .B2(new_n880), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n686), .A2(new_n281), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n913), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT57), .B1(new_n941), .B2(new_n518), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n684), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT59), .B(G148gat), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n935), .A2(new_n938), .A3(new_n945), .ZN(G1345gat));
  OAI21_X1  g745(.A(G155gat), .B1(new_n934), .B2(new_n711), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n711), .A2(G155gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n936), .B2(new_n948), .ZN(G1346gat));
  INV_X1    g748(.A(G162gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n950), .A3(new_n622), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n886), .A2(new_n621), .A3(new_n904), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n950), .B2(new_n952), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n746), .A2(new_n566), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n558), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n881), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(new_n386), .A3(new_n281), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n566), .B1(new_n877), .B2(new_n880), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n746), .A2(new_n579), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT124), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n735), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n958), .B1(new_n965), .B2(new_n386), .ZN(G1348gat));
  OAI21_X1  g765(.A(G176gat), .B1(new_n957), .B2(new_n685), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n684), .A2(new_n387), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G1349gat));
  NOR2_X1   g769(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n971));
  OAI21_X1  g770(.A(G183gat), .B1(new_n957), .B2(new_n711), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n959), .A2(new_n415), .A3(new_n667), .A4(new_n961), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g773(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n974), .B(new_n975), .ZN(G1350gat));
  NAND2_X1  g775(.A1(new_n621), .A2(new_n416), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n957), .B2(new_n622), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n980));
  OAI22_X1  g779(.A1(new_n968), .A2(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  NOR3_X1   g780(.A1(new_n703), .A2(new_n746), .A3(new_n519), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n959), .A2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n735), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n703), .A2(new_n955), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n986), .B1(new_n939), .B2(new_n942), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n280), .A2(G197gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(G1352gat));
  NOR3_X1   g789(.A1(new_n983), .A2(G204gat), .A3(new_n685), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  OAI21_X1  g793(.A(G204gat), .B1(new_n987), .B2(new_n685), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(G1353gat));
  OR3_X1    g795(.A1(new_n983), .A2(G211gat), .A3(new_n711), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n988), .A2(new_n667), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n998), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT63), .B1(new_n998), .B2(G211gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(G1354gat));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n622), .B1(new_n987), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1003), .B1(new_n1002), .B2(new_n987), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G218gat), .ZN(new_n1005));
  OR2_X1    g804(.A1(new_n622), .A2(G218gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n983), .B2(new_n1006), .ZN(G1355gat));
endmodule


