//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G217));
  OR4_X1    g027(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n440), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G125), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n466), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(G137), .A3(new_n470), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n470), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n472), .A2(new_n473), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n470), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT70), .Z(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n470), .C1(new_n472), .C2(new_n473), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n495), .A2(new_n506), .A3(new_n499), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n501), .A2(new_n504), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n520), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n519), .A2(G88), .B1(G651), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND2_X1  g108(.A1(new_n530), .A2(G51), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n519), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n534), .A2(new_n535), .A3(new_n537), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n510), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT73), .Z(new_n543));
  XOR2_X1   g118(.A(KEYINPUT74), .B(G90), .Z(new_n544));
  NAND2_X1  g119(.A1(new_n519), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n543), .B(new_n545), .C1(new_n546), .C2(new_n529), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n530), .A2(G43), .B1(G651), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n519), .A2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  AOI22_X1  g136(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n562), .B2(new_n510), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n525), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n516), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n572), .A2(new_n573), .A3(G53), .A4(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n519), .A2(G91), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(G299));
  AOI21_X1  g152(.A(G74), .B1(new_n522), .B2(new_n524), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT76), .B1(new_n578), .B2(new_n510), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n580), .B(G651), .C1(new_n517), .C2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n515), .A2(G49), .A3(G543), .A4(new_n516), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n572), .A2(G87), .A3(new_n517), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n530), .A2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n519), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n525), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n590), .A2(new_n591), .A3(G651), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n590), .B2(G651), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n586), .B(new_n587), .C1(new_n592), .C2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n519), .A2(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n530), .A2(G47), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n510), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n572), .A2(G92), .A3(new_n517), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n529), .A2(new_n603), .B1(new_n604), .B2(new_n510), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(G868), .B2(new_n608), .ZN(G284));
  OAI21_X1  g184(.A(new_n599), .B1(G868), .B2(new_n608), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NOR2_X1   g191(.A1(new_n555), .A2(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n608), .A2(new_n615), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n468), .A2(new_n479), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n486), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n488), .A2(G123), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2435), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2438), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  INV_X1    g213(.A(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(G1341), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2443), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n647), .A2(G14), .ZN(G401));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT81), .Z(new_n654));
  INV_X1    g229(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n649), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n655), .B(new_n656), .C1(new_n650), .C2(new_n651), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n655), .A2(new_n651), .A3(new_n649), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n631), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n669));
  INV_X1    g244(.A(new_n664), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  AOI22_X1  g246(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n664), .A3(new_n667), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n668), .C2(new_n669), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT83), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT84), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(G229));
  MUX2_X1   g259(.A(G24), .B(G290), .S(G16), .Z(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G1986), .Z(new_n686));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(KEYINPUT90), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G6), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n689), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n689), .A2(G23), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n579), .A2(new_n581), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n584), .A2(new_n583), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT89), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n582), .A2(new_n703), .A3(new_n583), .A4(new_n584), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n689), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT33), .B(G1976), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n694), .A2(new_n698), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n688), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n715));
  INV_X1    g290(.A(G95), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n470), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT86), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n486), .A2(G131), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n488), .A2(G119), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT87), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(new_n713), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n712), .B(new_n727), .C1(new_n711), .C2(new_n710), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT91), .Z(new_n729));
  AND2_X1   g304(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(G168), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G16), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n713), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n713), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT100), .B(KEYINPUT29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n713), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n713), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT99), .Z(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G2078), .ZN(new_n746));
  NOR2_X1   g321(.A1(G4), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n608), .B2(G16), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G1348), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n742), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n740), .A2(new_n741), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n745), .A2(G2078), .B1(G1348), .B2(new_n748), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT98), .B1(G5), .B2(G16), .ZN(new_n753));
  OR3_X1    g328(.A1(KEYINPUT98), .A2(G5), .A3(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(G301), .C2(new_n689), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n713), .B1(new_n758), .B2(G34), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(G34), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n483), .B2(new_n713), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  OR2_X1    g341(.A1(G29), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n486), .A2(G139), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n479), .A2(G103), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT94), .Z(new_n772));
  OAI211_X1 g347(.A(new_n768), .B(new_n770), .C1(new_n772), .C2(new_n470), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n713), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n765), .B1(new_n766), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n766), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT95), .Z(new_n777));
  NOR2_X1   g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT31), .B(G11), .Z(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n488), .A2(G129), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT97), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT26), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n486), .A2(G141), .B1(G105), .B2(new_n479), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n781), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT27), .B(G1996), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT93), .B(G2067), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n793));
  INV_X1    g368(.A(G26), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G29), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(G29), .ZN(new_n796));
  OR2_X1    g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT92), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n486), .A2(G140), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n488), .A2(G128), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(G29), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n795), .B1(new_n803), .B2(new_n793), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n791), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n555), .A2(new_n689), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n689), .B2(G19), .ZN(new_n807));
  INV_X1    g382(.A(G1341), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n734), .A2(new_n735), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n764), .A2(new_n757), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n808), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n804), .A2(new_n792), .ZN(new_n814));
  INV_X1    g389(.A(new_n630), .ZN(new_n815));
  INV_X1    g390(.A(G28), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT30), .ZN(new_n817));
  AOI21_X1  g392(.A(G29), .B1(new_n816), .B2(KEYINPUT30), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n815), .A2(G29), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n814), .B(new_n819), .C1(new_n755), .C2(new_n756), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n805), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT23), .B1(new_n612), .B2(new_n689), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n689), .A2(G20), .ZN(new_n823));
  MUX2_X1   g398(.A(KEYINPUT23), .B(new_n822), .S(new_n823), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G1956), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(G1956), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n779), .A2(new_n780), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n731), .A2(new_n732), .A3(new_n736), .A4(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n831), .A2(new_n529), .B1(new_n518), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n510), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  AND2_X1   g415(.A1(new_n835), .A2(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n554), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n555), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT39), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n608), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n840), .B1(new_n848), .B2(G860), .ZN(G145));
  INV_X1    g424(.A(G37), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n787), .B(new_n802), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n773), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n500), .A2(KEYINPUT102), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n495), .A2(new_n854), .A3(new_n499), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n504), .A2(new_n505), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n852), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n486), .A2(G142), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n488), .A2(G130), .ZN(new_n863));
  NOR2_X1   g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n623), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n722), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n493), .B(G160), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n630), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n868), .B(KEYINPUT103), .Z(new_n872));
  OAI211_X1 g447(.A(new_n869), .B(new_n871), .C1(new_n872), .C2(new_n861), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n861), .A2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n861), .A2(new_n872), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n850), .B(new_n873), .C1(new_n876), .C2(new_n871), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(G868), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n608), .B(G299), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n844), .B(new_n618), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G303), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n705), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n691), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n887), .B(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n887), .B1(new_n892), .B2(new_n891), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n884), .B2(new_n886), .ZN(new_n898));
  OAI22_X1  g473(.A1(new_n897), .A2(new_n898), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n879), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n841), .A2(G868), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(new_n900), .B2(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(new_n901), .A2(new_n904), .ZN(G331));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n844), .A2(G168), .ZN(new_n910));
  AOI21_X1  g485(.A(G286), .B1(new_n842), .B2(new_n843), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n910), .A2(G301), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(G301), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n881), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n880), .A3(new_n913), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT107), .A4(new_n880), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n890), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n912), .A2(new_n913), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n915), .B1(new_n922), .B2(new_n881), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n891), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n919), .A2(new_n890), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n927), .B2(new_n920), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n909), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n920), .A3(new_n921), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n920), .A2(new_n924), .ZN(new_n931));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n930), .C1(new_n931), .C2(new_n921), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(G397));
  AOI21_X1  g508(.A(G1384), .B1(new_n856), .B2(new_n858), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n935));
  XOR2_X1   g510(.A(KEYINPUT108), .B(G40), .Z(new_n936));
  AOI211_X1 g511(.A(new_n481), .B(new_n936), .C1(new_n471), .C2(new_n476), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n802), .B(G2067), .Z(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT110), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n941), .B2(new_n787), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n938), .A2(G1996), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n788), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n939), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n788), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT109), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(KEYINPUT109), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n722), .A2(new_n725), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n802), .A2(G2067), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n938), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n723), .A2(new_n726), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n939), .B1(new_n959), .B2(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n938), .A2(G1986), .A3(G290), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT48), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n947), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT125), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n967));
  AND2_X1   g542(.A1(G305), .A2(G1981), .ZN(new_n968));
  NOR2_X1   g543(.A1(G305), .A2(G1981), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT49), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n495), .A2(new_n854), .A3(new_n499), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n854), .B1(new_n495), .B2(new_n499), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n975), .B2(new_n857), .ZN(new_n976));
  INV_X1    g551(.A(new_n936), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT69), .B1(new_n475), .B2(G2105), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n465), .B(new_n470), .C1(new_n474), .C2(new_n466), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n482), .B(new_n977), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(G8), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n967), .B(new_n983), .C1(new_n968), .C2(new_n969), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n971), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n702), .B2(new_n704), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT52), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n981), .C2(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G288), .A2(new_n986), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n981), .A2(new_n987), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n985), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT45), .B(new_n972), .C1(new_n975), .C2(new_n857), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n937), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n508), .B2(new_n972), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G2078), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n508), .A2(new_n972), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n937), .A4(new_n999), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n980), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1012), .B(new_n972), .C1(new_n975), .C2(new_n857), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n859), .A2(KEYINPUT112), .A3(new_n1012), .A4(new_n972), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1009), .A2(new_n1010), .B1(new_n756), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(new_n937), .C1(new_n934), .C2(KEYINPUT45), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1010), .A2(G2078), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(G301), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n508), .A2(new_n1012), .A3(new_n972), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n937), .C1(new_n934), .C2(new_n1012), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G2090), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT113), .ZN(new_n1033));
  NAND3_X1  g608(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1030), .A2(new_n1035), .A3(new_n1031), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1029), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1017), .A2(G2090), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1037), .B(G8), .C1(new_n1025), .C2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n998), .A2(new_n1024), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(G286), .A2(G8), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1011), .A2(new_n1015), .A3(new_n757), .A4(new_n1016), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1020), .A2(new_n735), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1044), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT51), .B(G8), .C1(new_n1048), .C2(G286), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT62), .B(new_n1047), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n966), .B1(new_n1042), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1047), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1052), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT51), .B(new_n1043), .C1(new_n1048), .C2(G8), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n996), .B1(new_n990), .B2(new_n991), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1041), .A2(new_n985), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1008), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n980), .B1(new_n934), .B2(KEYINPUT45), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1007), .B1(new_n1063), .B2(new_n1006), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n697), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1028), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1037), .B1(new_n1067), .B2(G8), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1061), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1070), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1071), .A3(KEYINPUT125), .A4(new_n1024), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1054), .A2(new_n1059), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1017), .A2(new_n756), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(G301), .A3(new_n1075), .A4(new_n1023), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT54), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n475), .A2(G2105), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n1021), .C1(new_n934), .C2(KEYINPUT45), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n481), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n478), .A2(KEYINPUT122), .A3(new_n480), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1083), .A2(G40), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n999), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1078), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1022), .B1(new_n976), .B2(new_n1005), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(G40), .A3(new_n1083), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n934), .B2(KEYINPUT45), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1089), .A3(KEYINPUT123), .A4(new_n1079), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1018), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n998), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1074), .A2(new_n1091), .A3(G301), .A4(new_n1075), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT124), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1018), .A2(new_n1098), .A3(G301), .A4(new_n1091), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1074), .A2(new_n1075), .A3(new_n1023), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1956), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1027), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1063), .A2(new_n1006), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n575), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT118), .B1(new_n571), .B2(new_n574), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1115), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1116));
  OAI21_X1  g691(.A(G299), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT119), .B1(new_n1115), .B2(KEYINPUT57), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n612), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1109), .A2(new_n1121), .A3(KEYINPUT120), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT120), .B1(new_n1109), .B2(new_n1121), .ZN(new_n1123));
  INV_X1    g698(.A(new_n608), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n937), .A2(new_n934), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(G2067), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1017), .B2(new_n639), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1109), .A2(new_n1121), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1118), .A2(new_n612), .A3(new_n1119), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n612), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1136), .A2(new_n1107), .B1(new_n1105), .B2(new_n1027), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n608), .B(new_n1126), .C1(new_n639), .C2(new_n1017), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1106), .A2(new_n1108), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1129), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1006), .A2(new_n948), .A3(new_n937), .A4(new_n999), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n554), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1127), .A2(new_n1153), .A3(new_n608), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1146), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1131), .B1(new_n1143), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1095), .A2(new_n1104), .A3(new_n1156), .A4(new_n1058), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1060), .A2(new_n985), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n971), .A2(new_n984), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G288), .A2(G1976), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT116), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n969), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1158), .A2(new_n1041), .B1(new_n1162), .B2(new_n981), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1017), .A2(G2090), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1065), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1037), .B1(new_n1166), .B2(G8), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1164), .B1(new_n1167), .B2(new_n1158), .ZN(new_n1168));
  OAI21_X1  g743(.A(G8), .B1(new_n1025), .B2(new_n1040), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1038), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n998), .A2(KEYINPUT117), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1049), .A2(G286), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1172), .A2(new_n1041), .A3(KEYINPUT63), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n998), .A2(new_n1039), .A3(new_n1041), .A4(new_n1172), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1163), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1073), .A2(new_n1157), .A3(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(G1986), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n961), .B1(new_n939), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1179), .A2(KEYINPUT126), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT126), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n965), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(KEYINPUT127), .B(new_n965), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g763(.A1(G229), .A2(new_n463), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G401), .A2(G227), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1192), .A2(new_n877), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n927), .A2(new_n920), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1194), .A2(KEYINPUT43), .ZN(new_n1195));
  AOI211_X1 g769(.A(new_n1191), .B(new_n1193), .C1(new_n1195), .C2(new_n925), .ZN(G308));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n925), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n1197), .A2(new_n877), .A3(new_n1190), .A4(new_n1192), .ZN(G225));
endmodule


