

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752;

  XNOR2_X1 U375 ( .A(n535), .B(n534), .ZN(n751) );
  AND2_X1 U376 ( .A1(n536), .A2(n512), .ZN(n513) );
  XNOR2_X1 U377 ( .A(n462), .B(n461), .ZN(n470) );
  XNOR2_X1 U378 ( .A(n440), .B(n439), .ZN(n454) );
  XNOR2_X2 U379 ( .A(G143), .B(G128), .ZN(n440) );
  XNOR2_X2 U380 ( .A(n737), .B(G146), .ZN(n462) );
  BUF_X1 U381 ( .A(G128), .Z(n704) );
  AND2_X2 U382 ( .A1(n747), .A2(n520), .ZN(n521) );
  XNOR2_X2 U383 ( .A(n513), .B(KEYINPUT33), .ZN(n683) );
  XNOR2_X2 U384 ( .A(n579), .B(n578), .ZN(n600) );
  NAND2_X2 U385 ( .A1(n623), .A2(n510), .ZN(n525) );
  NOR2_X1 U386 ( .A1(n750), .A2(n748), .ZN(n584) );
  OR2_X1 U387 ( .A1(n533), .A2(n532), .ZN(n535) );
  NOR2_X1 U388 ( .A1(n385), .A2(n410), .ZN(n377) );
  XNOR2_X1 U389 ( .A(n390), .B(G119), .ZN(n468) );
  XNOR2_X1 U390 ( .A(KEYINPUT3), .B(G113), .ZN(n390) );
  NAND2_X1 U391 ( .A1(n616), .A2(n407), .ZN(n385) );
  OR2_X1 U392 ( .A1(n616), .A2(n383), .ZN(n382) );
  XNOR2_X2 U393 ( .A(n459), .B(n458), .ZN(n540) );
  XOR2_X1 U394 ( .A(G137), .B(G140), .Z(n479) );
  XNOR2_X1 U395 ( .A(G146), .B(G125), .ZN(n429) );
  NAND2_X1 U396 ( .A1(n382), .A2(n380), .ZN(n379) );
  NOR2_X1 U397 ( .A1(n381), .A2(n409), .ZN(n380) );
  INV_X1 U398 ( .A(KEYINPUT65), .ZN(n401) );
  XNOR2_X1 U399 ( .A(n400), .B(n399), .ZN(n726) );
  XNOR2_X1 U400 ( .A(KEYINPUT86), .B(G104), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n429), .B(n428), .ZN(n736) );
  XNOR2_X1 U402 ( .A(n427), .B(KEYINPUT10), .ZN(n428) );
  INV_X1 U403 ( .A(KEYINPUT67), .ZN(n427) );
  INV_X1 U404 ( .A(G107), .ZN(n361) );
  XNOR2_X1 U405 ( .A(n479), .B(n362), .ZN(n735) );
  INV_X1 U406 ( .A(KEYINPUT91), .ZN(n362) );
  XNOR2_X1 U407 ( .A(n726), .B(n461), .ZN(n457) );
  INV_X1 U408 ( .A(n379), .ZN(n374) );
  INV_X1 U409 ( .A(KEYINPUT98), .ZN(n365) );
  AND2_X1 U410 ( .A1(n529), .A2(n528), .ZN(n366) );
  XNOR2_X1 U411 ( .A(n444), .B(G478), .ZN(n445) );
  NOR2_X1 U412 ( .A1(n595), .A2(n594), .ZN(n598) );
  INV_X1 U413 ( .A(KEYINPUT78), .ZN(n369) );
  NAND2_X1 U414 ( .A1(n604), .A2(n555), .ZN(n370) );
  XNOR2_X1 U415 ( .A(n505), .B(KEYINPUT38), .ZN(n654) );
  NOR2_X1 U416 ( .A1(n669), .A2(n511), .ZN(n536) );
  NAND2_X1 U417 ( .A1(n407), .A2(n555), .ZN(n384) );
  INV_X1 U418 ( .A(G953), .ZN(n436) );
  INV_X1 U419 ( .A(G134), .ZN(n439) );
  XNOR2_X1 U420 ( .A(n432), .B(n431), .ZN(n608) );
  XNOR2_X1 U421 ( .A(n430), .B(n736), .ZN(n431) );
  XNOR2_X1 U422 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n396) );
  AND2_X1 U423 ( .A1(n604), .A2(n739), .ZN(n652) );
  NAND2_X1 U424 ( .A1(n374), .A2(n372), .ZN(n371) );
  NOR2_X1 U425 ( .A1(n373), .A2(KEYINPUT19), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n483), .B(n482), .ZN(n636) );
  XNOR2_X1 U427 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U428 ( .A(n457), .B(n359), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n735), .B(n360), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n456), .B(n361), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n612), .B(KEYINPUT85), .ZN(n650) );
  NAND2_X1 U432 ( .A1(n516), .A2(n560), .ZN(n519) );
  NAND2_X1 U433 ( .A1(n366), .A2(n364), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n508), .B(n365), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n460), .B(KEYINPUT99), .ZN(n489) );
  NAND2_X1 U436 ( .A1(n374), .A2(n385), .ZN(n355) );
  AND2_X1 U437 ( .A1(n382), .A2(n384), .ZN(n356) );
  OR2_X1 U438 ( .A1(n603), .A2(n602), .ZN(n357) );
  XNOR2_X1 U439 ( .A(n462), .B(n358), .ZN(n644) );
  XNOR2_X2 U440 ( .A(n363), .B(n509), .ZN(n623) );
  AND2_X4 U441 ( .A1(n627), .A2(n625), .ZN(n643) );
  XNOR2_X1 U442 ( .A(n370), .B(n369), .ZN(n368) );
  XNOR2_X2 U443 ( .A(n453), .B(KEYINPUT22), .ZN(n529) );
  NAND2_X2 U444 ( .A1(n367), .A2(n357), .ZN(n627) );
  NAND2_X1 U445 ( .A1(n368), .A2(n739), .ZN(n367) );
  NAND2_X2 U446 ( .A1(n375), .A2(n371), .ZN(n567) );
  INV_X1 U447 ( .A(n385), .ZN(n373) );
  AND2_X2 U448 ( .A1(n378), .A2(n376), .ZN(n375) );
  INV_X1 U449 ( .A(n377), .ZN(n376) );
  NAND2_X1 U450 ( .A1(n379), .A2(KEYINPUT19), .ZN(n378) );
  NAND2_X1 U451 ( .A1(n356), .A2(n385), .ZN(n505) );
  INV_X1 U452 ( .A(n384), .ZN(n381) );
  OR2_X1 U453 ( .A1(n407), .A2(n555), .ZN(n383) );
  BUF_X1 U454 ( .A(n436), .Z(n740) );
  AND2_X1 U455 ( .A1(n497), .A2(n663), .ZN(n386) );
  XOR2_X1 U456 ( .A(KEYINPUT7), .B(KEYINPUT94), .Z(n387) );
  XOR2_X1 U457 ( .A(n387), .B(n435), .Z(n388) );
  NOR2_X1 U458 ( .A1(n600), .A2(n599), .ZN(n389) );
  NOR2_X1 U459 ( .A1(G953), .A2(G237), .ZN(n463) );
  INV_X1 U460 ( .A(KEYINPUT19), .ZN(n410) );
  XNOR2_X1 U461 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U462 ( .A(KEYINPUT95), .ZN(n444) );
  XNOR2_X1 U463 ( .A(n488), .B(n487), .ZN(n663) );
  XNOR2_X1 U464 ( .A(n388), .B(n438), .ZN(n443) );
  XNOR2_X1 U465 ( .A(n446), .B(n445), .ZN(n544) );
  XNOR2_X1 U466 ( .A(n434), .B(n433), .ZN(n545) );
  XNOR2_X1 U467 ( .A(n443), .B(n442), .ZN(n640) );
  XNOR2_X1 U468 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n391) );
  XNOR2_X1 U469 ( .A(n468), .B(n391), .ZN(n393) );
  XNOR2_X1 U470 ( .A(G122), .B(G116), .ZN(n392) );
  XNOR2_X1 U471 ( .A(n392), .B(G107), .ZN(n441) );
  XNOR2_X1 U472 ( .A(n393), .B(n441), .ZN(n728) );
  NAND2_X1 U473 ( .A1(n436), .A2(G224), .ZN(n394) );
  XNOR2_X1 U474 ( .A(n394), .B(KEYINPUT4), .ZN(n395) );
  XNOR2_X1 U475 ( .A(n395), .B(n429), .ZN(n398) );
  XNOR2_X1 U476 ( .A(n440), .B(n396), .ZN(n397) );
  XNOR2_X1 U477 ( .A(n398), .B(n397), .ZN(n402) );
  INV_X1 U478 ( .A(G110), .ZN(n399) );
  XNOR2_X1 U479 ( .A(n401), .B(G101), .ZN(n461) );
  XNOR2_X1 U480 ( .A(n402), .B(n457), .ZN(n403) );
  XNOR2_X1 U481 ( .A(n728), .B(n403), .ZN(n616) );
  XNOR2_X1 U482 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  INV_X1 U483 ( .A(n603), .ZN(n555) );
  INV_X1 U484 ( .A(G902), .ZN(n484) );
  INV_X1 U485 ( .A(G237), .ZN(n404) );
  NAND2_X1 U486 ( .A1(n484), .A2(n404), .ZN(n408) );
  NAND2_X1 U487 ( .A1(n408), .A2(G210), .ZN(n406) );
  INV_X1 U488 ( .A(KEYINPUT87), .ZN(n405) );
  XNOR2_X1 U489 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U490 ( .A1(n408), .A2(G214), .ZN(n653) );
  INV_X1 U491 ( .A(n653), .ZN(n409) );
  NAND2_X1 U492 ( .A1(G234), .A2(G237), .ZN(n411) );
  XNOR2_X1 U493 ( .A(n411), .B(KEYINPUT14), .ZN(n415) );
  NAND2_X1 U494 ( .A1(n415), .A2(G902), .ZN(n412) );
  XOR2_X1 U495 ( .A(n412), .B(KEYINPUT89), .Z(n490) );
  INV_X1 U496 ( .A(n490), .ZN(n414) );
  XOR2_X1 U497 ( .A(G898), .B(KEYINPUT88), .Z(n723) );
  NAND2_X1 U498 ( .A1(G953), .A2(n723), .ZN(n729) );
  INV_X1 U499 ( .A(n729), .ZN(n413) );
  NAND2_X1 U500 ( .A1(n414), .A2(n413), .ZN(n417) );
  NAND2_X1 U501 ( .A1(G952), .A2(n415), .ZN(n681) );
  NOR2_X1 U502 ( .A1(n681), .A2(G953), .ZN(n495) );
  INV_X1 U503 ( .A(n495), .ZN(n416) );
  NAND2_X1 U504 ( .A1(n417), .A2(n416), .ZN(n418) );
  NAND2_X1 U505 ( .A1(n567), .A2(n418), .ZN(n419) );
  XNOR2_X2 U506 ( .A(n419), .B(KEYINPUT0), .ZN(n537) );
  XOR2_X1 U507 ( .A(KEYINPUT11), .B(KEYINPUT92), .Z(n421) );
  NAND2_X1 U508 ( .A1(G214), .A2(n463), .ZN(n420) );
  XNOR2_X1 U509 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U510 ( .A(n422), .B(G140), .Z(n432) );
  XOR2_X1 U511 ( .A(KEYINPUT12), .B(G104), .Z(n424) );
  XNOR2_X1 U512 ( .A(G143), .B(G131), .ZN(n423) );
  XNOR2_X1 U513 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U514 ( .A(G113), .B(G122), .Z(n425) );
  XNOR2_X1 U515 ( .A(n426), .B(n425), .ZN(n430) );
  NAND2_X1 U516 ( .A1(n608), .A2(n484), .ZN(n434) );
  XNOR2_X1 U517 ( .A(KEYINPUT13), .B(G475), .ZN(n433) );
  XNOR2_X1 U518 ( .A(KEYINPUT9), .B(KEYINPUT93), .ZN(n435) );
  NAND2_X1 U519 ( .A1(G234), .A2(n740), .ZN(n437) );
  XOR2_X1 U520 ( .A(KEYINPUT8), .B(n437), .Z(n477) );
  NAND2_X1 U521 ( .A1(G217), .A2(n477), .ZN(n438) );
  XNOR2_X1 U522 ( .A(n454), .B(n441), .ZN(n442) );
  NOR2_X1 U523 ( .A1(G902), .A2(n640), .ZN(n446) );
  NAND2_X1 U524 ( .A1(n545), .A2(n544), .ZN(n656) );
  INV_X1 U525 ( .A(n656), .ZN(n451) );
  NAND2_X1 U526 ( .A1(n603), .A2(G234), .ZN(n447) );
  XNOR2_X1 U527 ( .A(n447), .B(KEYINPUT20), .ZN(n485) );
  AND2_X1 U528 ( .A1(n485), .A2(G221), .ZN(n449) );
  INV_X1 U529 ( .A(KEYINPUT21), .ZN(n448) );
  XNOR2_X1 U530 ( .A(n449), .B(n448), .ZN(n662) );
  INV_X1 U531 ( .A(n662), .ZN(n450) );
  NAND2_X1 U532 ( .A1(n451), .A2(n450), .ZN(n452) );
  NOR2_X2 U533 ( .A1(n537), .A2(n452), .ZN(n453) );
  XNOR2_X1 U534 ( .A(KEYINPUT4), .B(G131), .ZN(n455) );
  XNOR2_X1 U535 ( .A(n455), .B(n454), .ZN(n737) );
  NAND2_X1 U536 ( .A1(G227), .A2(n740), .ZN(n456) );
  NAND2_X1 U537 ( .A1(n644), .A2(n484), .ZN(n459) );
  XNOR2_X1 U538 ( .A(KEYINPUT69), .B(G469), .ZN(n458) );
  XNOR2_X2 U539 ( .A(n540), .B(KEYINPUT1), .ZN(n511) );
  INV_X1 U540 ( .A(n511), .ZN(n501) );
  NAND2_X1 U541 ( .A1(n529), .A2(n511), .ZN(n460) );
  XOR2_X1 U542 ( .A(G116), .B(KEYINPUT5), .Z(n465) );
  NAND2_X1 U543 ( .A1(n463), .A2(G210), .ZN(n464) );
  XNOR2_X1 U544 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U545 ( .A(n466), .B(G137), .Z(n467) );
  XNOR2_X1 U546 ( .A(n470), .B(n469), .ZN(n630) );
  NAND2_X1 U547 ( .A1(n630), .A2(n484), .ZN(n473) );
  INV_X1 U548 ( .A(KEYINPUT72), .ZN(n471) );
  XNOR2_X1 U549 ( .A(n471), .B(G472), .ZN(n472) );
  XNOR2_X2 U550 ( .A(n473), .B(n472), .ZN(n497) );
  XOR2_X1 U551 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n475) );
  XNOR2_X1 U552 ( .A(n704), .B(KEYINPUT70), .ZN(n474) );
  XNOR2_X1 U553 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U554 ( .A(n736), .B(n476), .Z(n483) );
  NAND2_X1 U555 ( .A1(G221), .A2(n477), .ZN(n481) );
  XNOR2_X1 U556 ( .A(G110), .B(G119), .ZN(n478) );
  XNOR2_X1 U557 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U558 ( .A1(n636), .A2(n484), .ZN(n488) );
  NAND2_X1 U559 ( .A1(n485), .A2(G217), .ZN(n486) );
  XNOR2_X1 U560 ( .A(KEYINPUT25), .B(n486), .ZN(n487) );
  NAND2_X1 U561 ( .A1(n489), .A2(n386), .ZN(n510) );
  XNOR2_X1 U562 ( .A(n510), .B(G110), .ZN(G12) );
  OR2_X1 U563 ( .A1(n740), .A2(n490), .ZN(n491) );
  XNOR2_X1 U564 ( .A(KEYINPUT100), .B(n491), .ZN(n492) );
  NOR2_X1 U565 ( .A1(G900), .A2(n492), .ZN(n493) );
  XOR2_X1 U566 ( .A(KEYINPUT101), .B(n493), .Z(n494) );
  NOR2_X1 U567 ( .A1(n495), .A2(n494), .ZN(n574) );
  INV_X1 U568 ( .A(n663), .ZN(n531) );
  OR2_X1 U569 ( .A1(n531), .A2(n662), .ZN(n496) );
  NOR2_X1 U570 ( .A1(n574), .A2(n496), .ZN(n563) );
  XNOR2_X1 U571 ( .A(n497), .B(KEYINPUT6), .ZN(n512) );
  BUF_X1 U572 ( .A(n512), .Z(n507) );
  INV_X1 U573 ( .A(n545), .ZN(n498) );
  AND2_X1 U574 ( .A1(n498), .A2(n544), .ZN(n708) );
  AND2_X1 U575 ( .A1(n507), .A2(n708), .ZN(n499) );
  NAND2_X1 U576 ( .A1(n563), .A2(n499), .ZN(n500) );
  XNOR2_X1 U577 ( .A(KEYINPUT102), .B(n500), .ZN(n589) );
  NOR2_X1 U578 ( .A1(n589), .A2(n501), .ZN(n502) );
  NAND2_X1 U579 ( .A1(n653), .A2(n502), .ZN(n503) );
  XOR2_X1 U580 ( .A(KEYINPUT103), .B(n503), .Z(n504) );
  XNOR2_X1 U581 ( .A(n504), .B(KEYINPUT43), .ZN(n506) );
  AND2_X1 U582 ( .A1(n506), .A2(n505), .ZN(n601) );
  XOR2_X1 U583 ( .A(n601), .B(G140), .Z(G42) );
  INV_X1 U584 ( .A(n507), .ZN(n528) );
  XNOR2_X1 U585 ( .A(n511), .B(KEYINPUT83), .ZN(n591) );
  NAND2_X1 U586 ( .A1(n591), .A2(n663), .ZN(n508) );
  XNOR2_X1 U587 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n509) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT81), .ZN(n522) );
  NOR2_X1 U589 ( .A1(n662), .A2(n663), .ZN(n541) );
  INV_X1 U590 ( .A(n541), .ZN(n669) );
  XNOR2_X1 U591 ( .A(n537), .B(KEYINPUT90), .ZN(n542) );
  NOR2_X1 U592 ( .A1(n683), .A2(n542), .ZN(n515) );
  XOR2_X1 U593 ( .A(KEYINPUT34), .B(KEYINPUT75), .Z(n514) );
  XNOR2_X1 U594 ( .A(n515), .B(n514), .ZN(n516) );
  NOR2_X1 U595 ( .A1(n545), .A2(n544), .ZN(n560) );
  INV_X1 U596 ( .A(KEYINPUT74), .ZN(n517) );
  XNOR2_X1 U597 ( .A(n517), .B(KEYINPUT35), .ZN(n518) );
  XNOR2_X2 U598 ( .A(n519), .B(n518), .ZN(n747) );
  INV_X1 U599 ( .A(KEYINPUT44), .ZN(n520) );
  NAND2_X1 U600 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U601 ( .A(KEYINPUT71), .ZN(n523) );
  XNOR2_X1 U602 ( .A(n524), .B(n523), .ZN(n553) );
  INV_X1 U603 ( .A(n525), .ZN(n526) );
  NAND2_X1 U604 ( .A1(n747), .A2(n526), .ZN(n527) );
  NAND2_X1 U605 ( .A1(n527), .A2(KEYINPUT44), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U607 ( .A(n530), .B(KEYINPUT80), .ZN(n533) );
  NAND2_X1 U608 ( .A1(n511), .A2(n531), .ZN(n532) );
  INV_X1 U609 ( .A(KEYINPUT97), .ZN(n534) );
  INV_X1 U610 ( .A(n497), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n536), .A2(n556), .ZN(n674) );
  OR2_X1 U612 ( .A1(n674), .A2(n537), .ZN(n539) );
  INV_X1 U613 ( .A(KEYINPUT31), .ZN(n538) );
  XNOR2_X1 U614 ( .A(n539), .B(n538), .ZN(n714) );
  INV_X1 U615 ( .A(n540), .ZN(n565) );
  NAND2_X1 U616 ( .A1(n565), .A2(n541), .ZN(n573) );
  NOR2_X1 U617 ( .A1(n542), .A2(n573), .ZN(n543) );
  NAND2_X1 U618 ( .A1(n497), .A2(n543), .ZN(n696) );
  NAND2_X1 U619 ( .A1(n714), .A2(n696), .ZN(n548) );
  INV_X1 U620 ( .A(n544), .ZN(n546) );
  NAND2_X1 U621 ( .A1(n546), .A2(n545), .ZN(n715) );
  XNOR2_X1 U622 ( .A(KEYINPUT96), .B(n715), .ZN(n599) );
  INV_X1 U623 ( .A(n708), .ZN(n711) );
  NAND2_X1 U624 ( .A1(n599), .A2(n711), .ZN(n587) );
  INV_X1 U625 ( .A(n587), .ZN(n658) );
  XOR2_X1 U626 ( .A(KEYINPUT77), .B(n658), .Z(n571) );
  INV_X1 U627 ( .A(n571), .ZN(n547) );
  NAND2_X1 U628 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U629 ( .A1(n751), .A2(n549), .ZN(n550) );
  AND2_X1 U630 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U631 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X2 U632 ( .A(n554), .B(KEYINPUT45), .ZN(n604) );
  NAND2_X1 U633 ( .A1(n556), .A2(n653), .ZN(n557) );
  XNOR2_X1 U634 ( .A(n557), .B(KEYINPUT30), .ZN(n576) );
  OR2_X1 U635 ( .A1(n574), .A2(n576), .ZN(n558) );
  OR2_X1 U636 ( .A1(n573), .A2(n558), .ZN(n562) );
  INV_X1 U637 ( .A(n505), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n707) );
  AND2_X1 U640 ( .A1(n556), .A2(n563), .ZN(n564) );
  XNOR2_X1 U641 ( .A(KEYINPUT28), .B(n564), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n566), .A2(n565), .ZN(n582) );
  INV_X1 U643 ( .A(n567), .ZN(n568) );
  NOR2_X1 U644 ( .A1(n582), .A2(n568), .ZN(n709) );
  XOR2_X1 U645 ( .A(KEYINPUT47), .B(KEYINPUT66), .Z(n569) );
  NAND2_X1 U646 ( .A1(n709), .A2(n569), .ZN(n570) );
  NOR2_X1 U647 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U648 ( .A1(n707), .A2(n572), .ZN(n586) );
  OR2_X1 U649 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n577), .A2(n654), .ZN(n579) );
  INV_X1 U652 ( .A(KEYINPUT39), .ZN(n578) );
  NOR2_X1 U653 ( .A1(n600), .A2(n711), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n580), .B(KEYINPUT40), .ZN(n750) );
  NAND2_X1 U655 ( .A1(n654), .A2(n653), .ZN(n657) );
  NOR2_X1 U656 ( .A1(n656), .A2(n657), .ZN(n581) );
  XNOR2_X1 U657 ( .A(KEYINPUT41), .B(n581), .ZN(n684) );
  NOR2_X1 U658 ( .A1(n582), .A2(n684), .ZN(n583) );
  XNOR2_X1 U659 ( .A(KEYINPUT42), .B(n583), .ZN(n748) );
  XNOR2_X1 U660 ( .A(n584), .B(KEYINPUT46), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n709), .A2(n587), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n588), .A2(KEYINPUT47), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n589), .A2(n355), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n590), .B(KEYINPUT36), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n718) );
  NAND2_X1 U667 ( .A1(n593), .A2(n718), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n596) );
  XNOR2_X1 U669 ( .A(KEYINPUT79), .B(n596), .ZN(n597) );
  XNOR2_X1 U670 ( .A(n598), .B(n597), .ZN(n606) );
  NOR2_X1 U671 ( .A1(n601), .A2(n389), .ZN(n605) );
  INV_X1 U672 ( .A(KEYINPUT2), .ZN(n602) );
  AND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n739) );
  NAND2_X1 U674 ( .A1(n652), .A2(KEYINPUT2), .ZN(n625) );
  NAND2_X1 U675 ( .A1(n643), .A2(G475), .ZN(n610) );
  XNOR2_X1 U676 ( .A(KEYINPUT84), .B(KEYINPUT59), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(n613) );
  INV_X1 U679 ( .A(G952), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n611), .A2(G953), .ZN(n612) );
  NOR2_X2 U681 ( .A1(n613), .A2(n650), .ZN(n615) );
  XNOR2_X1 U682 ( .A(KEYINPUT64), .B(KEYINPUT60), .ZN(n614) );
  XNOR2_X1 U683 ( .A(n615), .B(n614), .ZN(G60) );
  NAND2_X1 U684 ( .A1(n643), .A2(G210), .ZN(n620) );
  XNOR2_X1 U685 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n617) );
  XOR2_X1 U686 ( .A(n617), .B(KEYINPUT55), .Z(n618) );
  XNOR2_X1 U687 ( .A(n616), .B(n618), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X2 U689 ( .A1(n621), .A2(n650), .ZN(n622) );
  XNOR2_X1 U690 ( .A(n622), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U691 ( .A(G119), .B(KEYINPUT126), .ZN(n624) );
  XNOR2_X1 U692 ( .A(n623), .B(n624), .ZN(G21) );
  AND2_X1 U693 ( .A1(n625), .A2(G472), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n632) );
  XNOR2_X1 U695 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT62), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U698 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U699 ( .A1(n633), .A2(n650), .ZN(n634) );
  XOR2_X1 U700 ( .A(n634), .B(KEYINPUT63), .Z(G57) );
  NAND2_X1 U701 ( .A1(n643), .A2(G217), .ZN(n638) );
  XNOR2_X1 U702 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U704 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n639), .A2(n650), .ZN(G66) );
  NAND2_X1 U706 ( .A1(n643), .A2(G478), .ZN(n641) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U708 ( .A1(n642), .A2(n650), .ZN(G63) );
  NAND2_X1 U709 ( .A1(n643), .A2(G469), .ZN(n649) );
  XOR2_X1 U710 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n646) );
  XNOR2_X1 U711 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n645) );
  XNOR2_X1 U712 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n644), .B(n647), .ZN(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n651), .A2(n650), .ZN(G54) );
  XNOR2_X1 U716 ( .A(n652), .B(KEYINPUT2), .ZN(n688) );
  NOR2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U718 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U720 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U721 ( .A1(n661), .A2(n683), .ZN(n679) );
  XOR2_X1 U722 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n665) );
  NAND2_X1 U723 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U724 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U725 ( .A(n666), .B(KEYINPUT114), .ZN(n667) );
  NOR2_X1 U726 ( .A1(n556), .A2(n667), .ZN(n668) );
  XNOR2_X1 U727 ( .A(n668), .B(KEYINPUT116), .ZN(n673) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n671) );
  NAND2_X1 U729 ( .A1(n511), .A2(n669), .ZN(n670) );
  XNOR2_X1 U730 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U733 ( .A(KEYINPUT51), .B(n676), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n677), .A2(n684), .ZN(n678) );
  NOR2_X1 U735 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n680), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U737 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U738 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U739 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n689), .B(KEYINPUT118), .ZN(n690) );
  NOR2_X1 U742 ( .A1(n690), .A2(G953), .ZN(n692) );
  XOR2_X1 U743 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n691) );
  XNOR2_X1 U744 ( .A(n692), .B(n691), .ZN(G75) );
  NOR2_X1 U745 ( .A1(n711), .A2(n696), .ZN(n694) );
  XNOR2_X1 U746 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n693) );
  XNOR2_X1 U747 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U748 ( .A(G104), .B(n695), .ZN(G6) );
  NOR2_X1 U749 ( .A1(n696), .A2(n715), .ZN(n700) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n698) );
  XNOR2_X1 U751 ( .A(G107), .B(KEYINPUT109), .ZN(n697) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(G9) );
  XOR2_X1 U754 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n703) );
  INV_X1 U755 ( .A(n715), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n709), .A2(n701), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n706) );
  XOR2_X1 U758 ( .A(n704), .B(KEYINPUT110), .Z(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(G30) );
  XOR2_X1 U760 ( .A(G143), .B(n707), .Z(G45) );
  NAND2_X1 U761 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U762 ( .A(G146), .B(n710), .ZN(G48) );
  NOR2_X1 U763 ( .A1(n711), .A2(n714), .ZN(n712) );
  XOR2_X1 U764 ( .A(KEYINPUT112), .B(n712), .Z(n713) );
  XNOR2_X1 U765 ( .A(G113), .B(n713), .ZN(G15) );
  NOR2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U767 ( .A(G116), .B(n716), .Z(G18) );
  XOR2_X1 U768 ( .A(G125), .B(KEYINPUT37), .Z(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(G27) );
  XNOR2_X1 U770 ( .A(G134), .B(n389), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n719), .B(KEYINPUT113), .ZN(G36) );
  INV_X1 U772 ( .A(n604), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n720), .A2(G953), .ZN(n725) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n721) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n721), .Z(n722) );
  NOR2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U777 ( .A1(n725), .A2(n724), .ZN(n732) );
  XOR2_X1 U778 ( .A(n726), .B(G101), .Z(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(n734) );
  XOR2_X1 U782 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n733) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(n738) );
  XOR2_X1 U785 ( .A(n738), .B(n737), .Z(n742) );
  XOR2_X1 U786 ( .A(n742), .B(n739), .Z(n741) );
  NAND2_X1 U787 ( .A1(n741), .A2(n740), .ZN(n746) );
  XNOR2_X1 U788 ( .A(G227), .B(n742), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(G900), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n744), .A2(G953), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n746), .A2(n745), .ZN(G72) );
  XNOR2_X1 U792 ( .A(n747), .B(G122), .ZN(G24) );
  XNOR2_X1 U793 ( .A(G137), .B(KEYINPUT127), .ZN(n749) );
  XNOR2_X1 U794 ( .A(n749), .B(n748), .ZN(G39) );
  XOR2_X1 U795 ( .A(G131), .B(n750), .Z(G33) );
  XNOR2_X1 U796 ( .A(G101), .B(KEYINPUT106), .ZN(n752) );
  XNOR2_X1 U797 ( .A(n752), .B(n751), .ZN(G3) );
endmodule

