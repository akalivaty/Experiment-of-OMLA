//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1221,
    new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT65), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .A3(G101), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G125), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n471), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n466), .A2(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n471), .B1(new_n464), .B2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n477), .C2(new_n478), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n471), .C1(new_n477), .C2(new_n478), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(new_n498), .A3(G138), .A4(new_n471), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n508), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n510), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n513), .A2(new_n512), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n509), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT70), .B1(new_n525), .B2(new_n530), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(new_n510), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT71), .B(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n516), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n538), .B(new_n540), .C1(new_n507), .C2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n507), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n510), .A2(new_n546), .B1(new_n516), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XNOR2_X1  g126(.A(KEYINPUT72), .B(KEYINPUT8), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT73), .ZN(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND3_X1  g131(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n527), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n539), .A2(G91), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n558), .A2(new_n562), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(G166), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n567), .B1(new_n508), .B2(new_n518), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(G303));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n507), .B1(new_n527), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n536), .B2(G49), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n516), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n516), .A2(new_n573), .A3(new_n574), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(G288));
  OAI211_X1 g153(.A(G48), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n516), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g156(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n513), .B2(new_n512), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n507), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n507), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n510), .A2(new_n594), .B1(new_n516), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n536), .A2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n527), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n505), .A2(new_n509), .A3(G92), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G321));
  NOR2_X1   g186(.A1(G299), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g188(.A(new_n612), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n615), .B2(G860), .ZN(G148));
  NOR2_X1   g191(.A1(new_n549), .A2(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n607), .A2(new_n608), .ZN(new_n618));
  INV_X1    g193(.A(new_n605), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G559), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT78), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n617), .B1(new_n622), .B2(G868), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n497), .A2(new_n469), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT12), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n497), .A2(new_n628), .A3(new_n469), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n466), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n486), .A2(G123), .ZN(new_n636));
  OR2_X1    g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT80), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n646), .B(new_n652), .Z(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n646), .B(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n655), .A2(G14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n666), .B1(new_n669), .B2(new_n663), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n663), .A3(new_n661), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n680), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n689), .A3(new_n684), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n682), .A2(new_n683), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n681), .A2(new_n685), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n682), .A3(new_n683), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(KEYINPUT83), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n686), .A2(new_n690), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G1981), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n696), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n679), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT84), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n691), .A2(KEYINPUT83), .A3(new_n695), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n709));
  OAI21_X1  g284(.A(G1981), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(G1986), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n704), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n704), .B2(new_n712), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n678), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n702), .A2(new_n703), .A3(new_n679), .ZN(new_n716));
  AOI21_X1  g291(.A(G1986), .B1(new_n710), .B2(new_n711), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n706), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n704), .A2(new_n707), .A3(new_n712), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n677), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n720), .ZN(G229));
  NOR2_X1   g296(.A1(G6), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n590), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n723), .B(new_n724), .Z(new_n725));
  NAND2_X1  g300(.A1(G288), .A2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G23), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT33), .B(G1976), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n727), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n727), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n725), .A2(new_n732), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n740));
  OAI21_X1  g315(.A(KEYINPUT85), .B1(new_n471), .B2(G107), .ZN(new_n741));
  OR2_X1    g316(.A1(G95), .A2(G2105), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n743), .B(G2104), .C1(new_n744), .C2(new_n742), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n486), .A2(G119), .ZN(new_n746));
  INV_X1    g321(.A(G131), .ZN(new_n747));
  INV_X1    g322(.A(new_n466), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G25), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT86), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n727), .A2(G24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n597), .B2(new_n727), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1986), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n752), .A2(new_n753), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n739), .A2(new_n740), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G21), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G168), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1966), .ZN(new_n767));
  INV_X1    g342(.A(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G27), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT94), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n496), .A2(new_n499), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n492), .A2(new_n493), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2078), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n768), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n466), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n486), .A2(G128), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT90), .B(G28), .Z(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n786), .B2(KEYINPUT30), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT30), .B2(new_n786), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n639), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(G29), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n727), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n549), .B2(new_n727), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n785), .B(new_n792), .C1(G1341), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n768), .A2(G32), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT89), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT26), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n466), .A2(G141), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n486), .A2(G129), .B1(G105), .B2(new_n469), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n768), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT27), .B(G1996), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  OR4_X1    g380(.A1(new_n767), .A2(new_n776), .A3(new_n795), .A4(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n497), .A2(G127), .ZN(new_n807));
  AND2_X1   g382(.A1(G115), .A2(G2104), .ZN(new_n808));
  OAI21_X1  g383(.A(G2105), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT25), .ZN(new_n810));
  NAND2_X1  g385(.A1(G103), .A2(G2104), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n471), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n466), .A2(G139), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G29), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G29), .B2(G33), .ZN(new_n817));
  INV_X1    g392(.A(G2072), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n819), .B(new_n820), .C1(G1341), .C2(new_n794), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n727), .A2(G20), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G299), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1956), .ZN(new_n826));
  INV_X1    g401(.A(G34), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(KEYINPUT24), .ZN(new_n828));
  AOI21_X1  g403(.A(G29), .B1(new_n827), .B2(KEYINPUT24), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(KEYINPUT87), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT87), .B2(new_n829), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT88), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n482), .B(KEYINPUT69), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n768), .ZN(new_n834));
  INV_X1    g409(.A(G2084), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(G5), .A2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT91), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G301), .B2(new_n727), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT92), .Z(new_n840));
  INV_X1    g415(.A(G1961), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n821), .A2(new_n826), .A3(new_n836), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n834), .A2(new_n835), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT93), .Z(new_n845));
  NOR2_X1   g420(.A1(G29), .A2(G35), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G162), .B2(G29), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G2090), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n727), .A2(G4), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n609), .B2(new_n727), .ZN(new_n853));
  INV_X1    g428(.A(G1348), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n851), .B(new_n855), .C1(new_n841), .C2(new_n840), .ZN(new_n856));
  NOR4_X1   g431(.A1(new_n806), .A2(new_n843), .A3(new_n845), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n763), .A2(new_n764), .A3(new_n857), .ZN(G150));
  INV_X1    g433(.A(G150), .ZN(G311));
  AOI22_X1  g434(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n507), .ZN(new_n861));
  INV_X1    g436(.A(G55), .ZN(new_n862));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n510), .A2(new_n862), .B1(new_n516), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT99), .B(G860), .Z(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n609), .A2(G559), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n549), .A2(new_n865), .ZN(new_n872));
  OAI22_X1  g447(.A1(new_n545), .A2(new_n548), .B1(new_n861), .B2(new_n864), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n871), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n866), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n868), .B1(new_n877), .B2(new_n879), .ZN(G145));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n466), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n486), .A2(G130), .ZN(new_n884));
  OR2_X1    g459(.A1(G106), .A2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n885), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n630), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n630), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n750), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n884), .A2(new_n886), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(new_n627), .A3(new_n629), .A4(new_n883), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n749), .A3(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n891), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n882), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n895), .ZN(new_n900));
  INV_X1    g475(.A(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT104), .A3(new_n896), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n809), .A2(new_n904), .A3(new_n814), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n802), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n904), .A3(new_n815), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n771), .A2(new_n911), .A3(new_n772), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(new_n783), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n783), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n909), .B1(new_n915), .B2(new_n914), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n899), .B(new_n903), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G160), .A2(new_n639), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n833), .A2(new_n791), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n920), .A2(new_n921), .A3(G162), .ZN(new_n922));
  AOI21_X1  g497(.A(G162), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n897), .A2(new_n882), .A3(new_n898), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n914), .A2(new_n915), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n906), .A2(new_n908), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n928), .A3(new_n916), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n919), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n924), .B1(new_n919), .B2(new_n929), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n881), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n919), .A2(new_n929), .ZN(new_n935));
  INV_X1    g510(.A(new_n924), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .A3(new_n931), .A4(new_n930), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(G395));
  INV_X1    g516(.A(G288), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n590), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G166), .B(new_n597), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n588), .A2(G288), .A3(new_n589), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(KEYINPUT111), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n872), .A2(new_n873), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT107), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n622), .B(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n620), .A2(new_n956), .A3(G299), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT9), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n557), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n562), .A2(new_n563), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n558), .A2(KEYINPUT108), .A3(new_n562), .A4(new_n563), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n609), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(KEYINPUT109), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(KEYINPUT109), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n955), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT110), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n957), .A2(new_n963), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n957), .B2(new_n963), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n968), .B(KEYINPUT110), .C1(new_n955), .C2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n952), .A2(new_n969), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n952), .B1(new_n974), .B2(new_n969), .ZN(new_n976));
  OAI21_X1  g551(.A(G868), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n865), .A2(G868), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(G295));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n978), .ZN(G331));
  NAND2_X1  g555(.A1(G168), .A2(G171), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n533), .A2(G301), .A3(new_n534), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n874), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n533), .A2(G301), .A3(new_n534), .ZN(new_n984));
  AOI21_X1  g559(.A(G301), .B1(new_n533), .B2(new_n534), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n953), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n971), .B2(new_n972), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n946), .A2(new_n947), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n964), .A2(new_n983), .A3(new_n986), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n931), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n988), .B2(new_n990), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT112), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n983), .B(new_n986), .C1(new_n965), .C2(new_n966), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n973), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n987), .B1(new_n971), .B2(KEYINPUT113), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n996), .B(new_n948), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n931), .A4(new_n991), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(KEYINPUT43), .C1(new_n992), .C2(new_n993), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n995), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1001), .B1(new_n992), .B2(new_n993), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n931), .A3(new_n991), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n1001), .ZN(new_n1008));
  MUX2_X1   g583(.A(new_n1005), .B(new_n1008), .S(KEYINPUT44), .Z(G397));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  INV_X1    g585(.A(G40), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n476), .A2(new_n1011), .A3(new_n481), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n771), .B2(new_n772), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n572), .B(G1976), .C1(new_n576), .C2(new_n577), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G1981), .B1(new_n581), .B2(new_n586), .ZN(new_n1022));
  INV_X1    g597(.A(G61), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n503), .B2(new_n504), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G73), .A2(G543), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT76), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G651), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n505), .A2(new_n509), .A3(G86), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n701), .A3(new_n1031), .A4(new_n579), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1022), .A2(KEYINPUT117), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(G1981), .C1(new_n581), .C2(new_n586), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(KEYINPUT119), .A3(KEYINPUT49), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1014), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1033), .A2(new_n1043), .A3(new_n1035), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1033), .A2(KEYINPUT118), .A3(new_n1043), .A4(new_n1035), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1021), .B1(new_n1041), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n479), .A2(new_n480), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G2105), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(G40), .A3(new_n467), .A4(new_n475), .ZN(new_n1052));
  INV_X1    g627(.A(G1384), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n773), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n910), .A2(KEYINPUT45), .A3(new_n1053), .A4(new_n912), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1971), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1052), .B1(new_n1013), .B2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1061), .A3(new_n850), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n566), .A2(G8), .A3(new_n568), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n566), .A2(G8), .A3(new_n568), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1013), .B2(new_n1060), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT115), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n835), .A3(new_n1061), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1010), .B(G286), .C1(new_n1077), .C2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1076), .A2(new_n850), .A3(new_n1061), .ZN(new_n1083));
  OAI211_X1 g658(.A(G8), .B(new_n1070), .C1(new_n1083), .C2(new_n1058), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1049), .A2(new_n1072), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n736), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1076), .A2(new_n850), .A3(new_n1061), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1010), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1091), .B2(new_n1070), .ZN(new_n1092));
  OAI21_X1  g667(.A(G8), .B1(new_n1083), .B2(new_n1058), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1071), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1092), .A2(new_n1094), .A3(new_n1049), .A4(new_n1082), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n942), .A2(new_n1018), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1041), .B2(new_n1048), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1032), .B(KEYINPUT120), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1014), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1049), .A2(new_n1091), .A3(new_n1070), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1100), .A2(KEYINPUT121), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT121), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1096), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT122), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1077), .A2(G168), .A3(new_n1081), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT51), .B1(new_n1106), .B2(G8), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1110), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(G8), .A3(G286), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1112), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n1120), .B2(new_n1116), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1088), .B2(G2078), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1076), .A2(new_n1061), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n841), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1122), .A2(G2078), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1056), .B(new_n1127), .C1(new_n1055), .C2(new_n1054), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1049), .A2(new_n1084), .A3(new_n1072), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1129), .A2(new_n1130), .A3(G301), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1119), .A2(new_n1121), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1056), .A2(new_n1057), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT123), .ZN(new_n1140));
  XOR2_X1   g715(.A(G299), .B(KEYINPUT57), .Z(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1124), .A2(new_n854), .ZN(new_n1145));
  INV_X1    g720(.A(G2067), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1012), .A2(new_n1013), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n620), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1140), .A2(new_n1143), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1141), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1141), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1144), .A2(KEYINPUT61), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT58), .B(G1341), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1054), .B2(new_n1052), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT124), .B(G1996), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1088), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(KEYINPUT59), .A3(new_n549), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n549), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1153), .A2(new_n1154), .A3(new_n1159), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n609), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n620), .A4(new_n1147), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(new_n1165), .B2(new_n1164), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1149), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1170));
  XNOR2_X1  g745(.A(G301), .B(KEYINPUT54), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n910), .A2(new_n1053), .A3(new_n912), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1055), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1173), .A2(new_n1012), .A3(new_n1057), .A4(new_n1127), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1126), .B2(new_n1174), .ZN(new_n1175));
  AND4_X1   g750(.A1(new_n1128), .A2(new_n1123), .A3(new_n1125), .A4(new_n1171), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n1130), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1169), .A2(new_n1170), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1096), .B(new_n1180), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1105), .A2(new_n1132), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT114), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n1173), .B2(new_n1052), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1172), .A2(KEYINPUT114), .A3(new_n1055), .A4(new_n1012), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(G1996), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n907), .B(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n783), .B(new_n1146), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n750), .A2(new_n753), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n750), .A2(new_n753), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n597), .B(new_n679), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1186), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1182), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1184), .A2(new_n1187), .A3(new_n1185), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT46), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n802), .A2(new_n1189), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1186), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1197), .A2(KEYINPUT47), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT47), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1202));
  OR3_X1    g777(.A1(new_n1201), .A2(KEYINPUT126), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT126), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1186), .A2(new_n679), .A3(new_n597), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1205), .A2(KEYINPUT48), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1205), .A2(KEYINPUT48), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1208), .A2(new_n1190), .B1(G2067), .B2(new_n783), .ZN(new_n1209));
  AOI22_X1  g784(.A1(new_n1206), .A2(new_n1207), .B1(new_n1186), .B2(new_n1209), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1203), .A2(new_n1204), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g787(.A1(new_n659), .A2(new_n462), .A3(G227), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n715), .A2(new_n720), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1215), .B1(new_n934), .B2(new_n938), .ZN(new_n1216));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n1216), .A2(new_n1217), .A3(new_n1005), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n1217), .B1(new_n1216), .B2(new_n1005), .ZN(new_n1219));
  NOR2_X1   g793(.A1(new_n1218), .A2(new_n1219), .ZN(G308));
  NAND2_X1  g794(.A1(new_n1216), .A2(new_n1005), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1221), .A2(KEYINPUT127), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n1216), .A2(new_n1217), .A3(new_n1005), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1223), .ZN(G225));
endmodule


