

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U550 ( .A1(n707), .A2(n631), .ZN(n653) );
  INV_X2 U551 ( .A(n706), .ZN(n631) );
  NOR2_X1 U552 ( .A1(n740), .A2(n739), .ZN(n742) );
  OR2_X1 U553 ( .A1(n636), .A2(n635), .ZN(n641) );
  AND2_X1 U554 ( .A1(n670), .A2(n667), .ZN(n668) );
  AND2_X1 U555 ( .A1(n735), .A2(n729), .ZN(n516) );
  NOR2_X1 U556 ( .A1(n991), .A2(n624), .ZN(n627) );
  INV_X1 U557 ( .A(KEYINPUT100), .ZN(n639) );
  AND2_X1 U558 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U559 ( .A(n679), .B(KEYINPUT102), .ZN(n680) );
  XNOR2_X1 U560 ( .A(n687), .B(KEYINPUT104), .ZN(n688) );
  NOR2_X1 U561 ( .A1(n688), .A2(n733), .ZN(n689) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  INV_X1 U564 ( .A(KEYINPUT105), .ZN(n741) );
  INV_X1 U565 ( .A(KEYINPUT14), .ZN(n608) );
  INV_X1 U566 ( .A(G2104), .ZN(n528) );
  XNOR2_X1 U567 ( .A(n609), .B(n608), .ZN(n615) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n539), .Z(n784) );
  NOR2_X1 U569 ( .A1(G651), .A2(n575), .ZN(n787) );
  NAND2_X1 U570 ( .A1(n528), .A2(G2105), .ZN(n517) );
  XNOR2_X2 U571 ( .A(n517), .B(KEYINPUT65), .ZN(n886) );
  NAND2_X1 U572 ( .A1(G125), .A2(n886), .ZN(n518) );
  XNOR2_X1 U573 ( .A(n518), .B(KEYINPUT66), .ZN(n527) );
  INV_X1 U574 ( .A(KEYINPUT67), .ZN(n522) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT17), .ZN(n532) );
  INV_X1 U576 ( .A(G137), .ZN(n520) );
  OR2_X1 U577 ( .A1(n532), .A2(n520), .ZN(n521) );
  XNOR2_X1 U578 ( .A(n522), .B(n521), .ZN(n524) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U580 ( .A1(n888), .A2(G113), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U582 ( .A(KEYINPUT68), .B(n525), .Z(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n531) );
  NOR2_X1 U584 ( .A1(G2105), .A2(n528), .ZN(n882) );
  NAND2_X1 U585 ( .A1(G101), .A2(n882), .ZN(n529) );
  XNOR2_X1 U586 ( .A(KEYINPUT23), .B(n529), .ZN(n530) );
  NOR2_X2 U587 ( .A1(n531), .A2(n530), .ZN(G160) );
  NAND2_X1 U588 ( .A1(G102), .A2(n882), .ZN(n534) );
  INV_X1 U589 ( .A(n532), .ZN(n883) );
  NAND2_X1 U590 ( .A1(n883), .A2(G138), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G114), .A2(n888), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G126), .A2(n886), .ZN(n535) );
  NAND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n538), .A2(n537), .ZN(G164) );
  XOR2_X1 U596 ( .A(G651), .B(KEYINPUT70), .Z(n541) );
  NOR2_X1 U597 ( .A1(G543), .A2(n541), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G65), .A2(n784), .ZN(n543) );
  XNOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U600 ( .A(n540), .B(KEYINPUT69), .ZN(n575) );
  NOR2_X1 U601 ( .A1(n575), .A2(n541), .ZN(n791) );
  NAND2_X1 U602 ( .A1(G78), .A2(n791), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n546) );
  NOR2_X1 U604 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U605 ( .A1(n783), .A2(G91), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT74), .B(n544), .Z(n545) );
  NOR2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n787), .A2(G53), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U610 ( .A1(n787), .A2(G52), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G64), .A2(n784), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U613 ( .A(KEYINPUT72), .B(n551), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G90), .A2(n783), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G77), .A2(n791), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G171) );
  NAND2_X1 U619 ( .A1(n783), .A2(G89), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G76), .A2(n791), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n560), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U624 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n787), .A2(G51), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G63), .A2(n784), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G88), .A2(n783), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT84), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G62), .A2(n784), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n787), .A2(G50), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G75), .A2(n791), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(G166) );
  INV_X1 U640 ( .A(G166), .ZN(G303) );
  NAND2_X1 U641 ( .A1(G87), .A2(n575), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G49), .A2(n787), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n784), .A2(n578), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT81), .B(n579), .Z(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT82), .ZN(G288) );
  NAND2_X1 U649 ( .A1(n783), .A2(G86), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G61), .A2(n784), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G73), .A2(n791), .ZN(n585) );
  XOR2_X1 U653 ( .A(KEYINPUT2), .B(n585), .Z(n586) );
  NOR2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U655 ( .A(KEYINPUT83), .B(n588), .Z(n590) );
  NAND2_X1 U656 ( .A1(n787), .A2(G48), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(G305) );
  NAND2_X1 U658 ( .A1(G85), .A2(n783), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G72), .A2(n791), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G60), .A2(n784), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n787), .A2(G47), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(G290) );
  NAND2_X1 U666 ( .A1(G160), .A2(G40), .ZN(n706) );
  INV_X1 U667 ( .A(n653), .ZN(n646) );
  AND2_X1 U668 ( .A1(n646), .A2(G2067), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT99), .ZN(n600) );
  INV_X1 U670 ( .A(n646), .ZN(n671) );
  NAND2_X1 U671 ( .A1(n671), .A2(G1348), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n626) );
  NAND2_X1 U673 ( .A1(n783), .A2(G92), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G66), .A2(n784), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n787), .A2(G54), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G79), .A2(n791), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT15), .B(n607), .Z(n977) );
  NAND2_X1 U681 ( .A1(n784), .A2(G56), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n783), .A2(G81), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G68), .A2(n791), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U686 ( .A(KEYINPUT13), .B(n613), .Z(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n787), .A2(G43), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n991) );
  AND2_X1 U690 ( .A1(G160), .A2(G40), .ZN(n619) );
  AND2_X1 U691 ( .A1(G1996), .A2(n707), .ZN(n618) );
  AND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n653), .A2(G1341), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n977), .A2(n627), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n629) );
  OR2_X1 U699 ( .A1(n977), .A2(n627), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n638) );
  NAND2_X1 U701 ( .A1(n653), .A2(G1956), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(KEYINPUT97), .ZN(n636) );
  XOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n634) );
  AND2_X1 U704 ( .A1(n707), .A2(G2072), .ZN(n632) );
  AND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n635) );
  OR2_X1 U707 ( .A1(G299), .A2(n641), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n644) );
  NAND2_X1 U710 ( .A1(G299), .A2(n641), .ZN(n642) );
  XOR2_X1 U711 ( .A(KEYINPUT28), .B(n642), .Z(n643) );
  NOR2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n645), .B(KEYINPUT29), .ZN(n651) );
  XOR2_X1 U714 ( .A(G2078), .B(KEYINPUT25), .Z(n953) );
  NOR2_X1 U715 ( .A1(n953), .A2(n671), .ZN(n648) );
  XNOR2_X1 U716 ( .A(G1961), .B(KEYINPUT94), .ZN(n998) );
  NOR2_X1 U717 ( .A1(n646), .A2(n998), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT95), .B(n649), .ZN(n652) );
  NAND2_X1 U720 ( .A1(G171), .A2(n652), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n661) );
  NOR2_X1 U722 ( .A1(G171), .A2(n652), .ZN(n658) );
  NAND2_X1 U723 ( .A1(G8), .A2(n653), .ZN(n733) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n733), .ZN(n664) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n653), .ZN(n662) );
  NOR2_X1 U726 ( .A1(n664), .A2(n662), .ZN(n654) );
  NAND2_X1 U727 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U729 ( .A1(G168), .A2(n656), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U731 ( .A(KEYINPUT31), .B(n659), .Z(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n670) );
  NAND2_X1 U733 ( .A1(G8), .A2(n662), .ZN(n663) );
  XOR2_X1 U734 ( .A(KEYINPUT93), .B(n663), .Z(n666) );
  INV_X1 U735 ( .A(n664), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT101), .B(n668), .ZN(n683) );
  AND2_X1 U737 ( .A1(G286), .A2(G8), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n678) );
  INV_X1 U739 ( .A(G8), .ZN(n676) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n733), .ZN(n673) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n671), .ZN(n672) );
  NOR2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n674), .A2(G303), .ZN(n675) );
  OR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n681) );
  INV_X1 U746 ( .A(KEYINPUT32), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n722) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n732) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n732), .A2(n684), .ZN(n984) );
  NAND2_X1 U752 ( .A1(n722), .A2(n984), .ZN(n686) );
  NAND2_X1 U753 ( .A1(G288), .A2(G1976), .ZN(n685) );
  XOR2_X1 U754 ( .A(KEYINPUT103), .B(n685), .Z(n988) );
  NAND2_X1 U755 ( .A1(n686), .A2(n988), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n689), .B(KEYINPUT64), .ZN(n731) );
  NAND2_X1 U757 ( .A1(G117), .A2(n888), .ZN(n691) );
  NAND2_X1 U758 ( .A1(G129), .A2(n886), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n882), .A2(G105), .ZN(n692) );
  XOR2_X1 U761 ( .A(KEYINPUT38), .B(n692), .Z(n693) );
  NOR2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n883), .A2(G141), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n862) );
  NAND2_X1 U765 ( .A1(G1996), .A2(n862), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(KEYINPUT91), .ZN(n705) );
  INV_X1 U767 ( .A(G1991), .ZN(n949) );
  NAND2_X1 U768 ( .A1(G95), .A2(n882), .ZN(n699) );
  NAND2_X1 U769 ( .A1(G131), .A2(n883), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G107), .A2(n888), .ZN(n701) );
  NAND2_X1 U772 ( .A1(G119), .A2(n886), .ZN(n700) );
  NAND2_X1 U773 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n863) );
  NOR2_X1 U775 ( .A1(n949), .A2(n863), .ZN(n704) );
  NOR2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n926) );
  NOR2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n755) );
  INV_X1 U778 ( .A(n755), .ZN(n708) );
  NOR2_X1 U779 ( .A1(n926), .A2(n708), .ZN(n747) );
  INV_X1 U780 ( .A(n747), .ZN(n719) );
  XNOR2_X1 U781 ( .A(G2067), .B(KEYINPUT37), .ZN(n752) );
  NAND2_X1 U782 ( .A1(G116), .A2(n888), .ZN(n710) );
  NAND2_X1 U783 ( .A1(G128), .A2(n886), .ZN(n709) );
  NAND2_X1 U784 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U785 ( .A(n711), .B(KEYINPUT35), .ZN(n716) );
  NAND2_X1 U786 ( .A1(G104), .A2(n882), .ZN(n713) );
  NAND2_X1 U787 ( .A1(G140), .A2(n883), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U789 ( .A(KEYINPUT34), .B(n714), .Z(n715) );
  NAND2_X1 U790 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U791 ( .A(n717), .B(KEYINPUT36), .Z(n864) );
  OR2_X1 U792 ( .A1(n752), .A2(n864), .ZN(n718) );
  XOR2_X1 U793 ( .A(KEYINPUT90), .B(n718), .Z(n940) );
  NAND2_X1 U794 ( .A1(n755), .A2(n940), .ZN(n750) );
  AND2_X1 U795 ( .A1(n719), .A2(n750), .ZN(n735) );
  NOR2_X1 U796 ( .A1(G2090), .A2(G303), .ZN(n720) );
  NAND2_X1 U797 ( .A1(G8), .A2(n720), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U799 ( .A1(n723), .A2(n733), .ZN(n728) );
  NOR2_X1 U800 ( .A1(G1981), .A2(G305), .ZN(n724) );
  XOR2_X1 U801 ( .A(n724), .B(KEYINPUT24), .Z(n725) );
  NOR2_X1 U802 ( .A1(n733), .A2(n725), .ZN(n726) );
  XOR2_X1 U803 ( .A(n726), .B(KEYINPUT92), .Z(n727) );
  NAND2_X1 U804 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U805 ( .A1(KEYINPUT33), .A2(n516), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n740) );
  NAND2_X1 U807 ( .A1(n732), .A2(KEYINPUT33), .ZN(n734) );
  NOR2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n737) );
  XOR2_X1 U809 ( .A(G1981), .B(G305), .Z(n974) );
  NAND2_X1 U810 ( .A1(n974), .A2(n735), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U812 ( .A1(n516), .A2(n738), .ZN(n739) );
  XNOR2_X1 U813 ( .A(n742), .B(n741), .ZN(n744) );
  XNOR2_X1 U814 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U815 ( .A1(n981), .A2(n755), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n758) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n862), .ZN(n934) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n745) );
  AND2_X1 U819 ( .A1(n949), .A2(n863), .ZN(n924) );
  NOR2_X1 U820 ( .A1(n745), .A2(n924), .ZN(n746) );
  NOR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n934), .A2(n748), .ZN(n749) );
  XNOR2_X1 U823 ( .A(n749), .B(KEYINPUT39), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n864), .A2(n752), .ZN(n922) );
  NAND2_X1 U826 ( .A1(n753), .A2(n922), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U828 ( .A(KEYINPUT106), .B(n756), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U831 ( .A1(G99), .A2(n882), .ZN(n761) );
  NAND2_X1 U832 ( .A1(G111), .A2(n888), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n886), .A2(G123), .ZN(n762) );
  XOR2_X1 U835 ( .A(KEYINPUT18), .B(n762), .Z(n763) );
  NOR2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n883), .A2(G135), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n766), .A2(n765), .ZN(n921) );
  XNOR2_X1 U839 ( .A(G2096), .B(n921), .ZN(n767) );
  OR2_X1 U840 ( .A1(G2100), .A2(n767), .ZN(G156) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  NAND2_X1 U843 ( .A1(G94), .A2(G452), .ZN(n768) );
  XNOR2_X1 U844 ( .A(n768), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n769) );
  XNOR2_X1 U846 ( .A(n769), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U847 ( .A(G223), .ZN(n827) );
  NAND2_X1 U848 ( .A1(n827), .A2(G567), .ZN(n770) );
  XOR2_X1 U849 ( .A(KEYINPUT11), .B(n770), .Z(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n795) );
  OR2_X1 U851 ( .A1(n991), .A2(n795), .ZN(G153) );
  INV_X1 U852 ( .A(G171), .ZN(G301) );
  INV_X1 U853 ( .A(n977), .ZN(n778) );
  NOR2_X1 U854 ( .A1(G868), .A2(n778), .ZN(n772) );
  INV_X1 U855 ( .A(G868), .ZN(n809) );
  NOR2_X1 U856 ( .A1(n809), .A2(G301), .ZN(n771) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U858 ( .A(KEYINPUT76), .B(n773), .ZN(G284) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n775) );
  NOR2_X1 U860 ( .A1(G286), .A2(n809), .ZN(n774) );
  NOR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n795), .A2(G559), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n776), .A2(n977), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(n778), .A2(n809), .ZN(n779) );
  XOR2_X1 U866 ( .A(KEYINPUT78), .B(n779), .Z(n780) );
  NOR2_X1 U867 ( .A1(G559), .A2(n780), .ZN(n782) );
  NOR2_X1 U868 ( .A1(G868), .A2(n991), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U870 ( .A1(n783), .A2(G93), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G67), .A2(n784), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U873 ( .A1(n787), .A2(G55), .ZN(n788) );
  XOR2_X1 U874 ( .A(KEYINPUT80), .B(n788), .Z(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G80), .A2(n791), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n793), .A2(n792), .ZN(n808) );
  NAND2_X1 U878 ( .A1(G559), .A2(n977), .ZN(n794) );
  XOR2_X1 U879 ( .A(n991), .B(n794), .Z(n806) );
  NAND2_X1 U880 ( .A1(n795), .A2(n806), .ZN(n796) );
  XNOR2_X1 U881 ( .A(n796), .B(KEYINPUT79), .ZN(n797) );
  XOR2_X1 U882 ( .A(n808), .B(n797), .Z(G145) );
  XOR2_X1 U883 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n799) );
  XNOR2_X1 U884 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n798) );
  XNOR2_X1 U885 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U886 ( .A(G166), .B(n800), .ZN(n802) );
  XNOR2_X1 U887 ( .A(G290), .B(G288), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n802), .B(n801), .ZN(n803) );
  XOR2_X1 U889 ( .A(n808), .B(n803), .Z(n805) );
  XOR2_X1 U890 ( .A(G305), .B(G299), .Z(n804) );
  XNOR2_X1 U891 ( .A(n805), .B(n804), .ZN(n899) );
  XNOR2_X1 U892 ( .A(n806), .B(n899), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n807), .A2(G868), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U895 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U901 ( .A(KEYINPUT75), .B(G57), .ZN(G237) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U903 ( .A1(G108), .A2(G120), .ZN(n816) );
  NOR2_X1 U904 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G69), .A2(n817), .ZN(n832) );
  NAND2_X1 U906 ( .A1(G567), .A2(n832), .ZN(n822) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n818) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n818), .Z(n819) );
  NOR2_X1 U909 ( .A1(G218), .A2(n819), .ZN(n820) );
  NAND2_X1 U910 ( .A1(G96), .A2(n820), .ZN(n833) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n833), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT88), .B(n823), .Z(G319) );
  INV_X1 U914 ( .A(G319), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G661), .A2(G483), .ZN(n824) );
  NOR2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT89), .B(n826), .Z(n830) );
  NAND2_X1 U918 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U924 ( .A(KEYINPUT109), .B(n831), .Z(G188) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G108), .ZN(G238) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n835) );
  XNOR2_X1 U933 ( .A(KEYINPUT110), .B(G2096), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n836), .B(KEYINPUT42), .Z(n838) );
  XNOR2_X1 U936 ( .A(G2072), .B(G2067), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U938 ( .A(G2100), .B(G2084), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2090), .B(G2078), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2678), .B(KEYINPUT111), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U944 ( .A(G1966), .B(G1956), .Z(n846) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1961), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U948 ( .A(G1976), .B(G1971), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1991), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1981), .B(G1996), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G100), .A2(n882), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G136), .A2(n883), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G124), .A2(n886), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G112), .A2(n888), .ZN(n857) );
  XOR2_X1 U960 ( .A(KEYINPUT113), .B(n857), .Z(n858) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n867) );
  XNOR2_X1 U966 ( .A(G164), .B(KEYINPUT115), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(n869), .B(n868), .Z(n881) );
  NAND2_X1 U969 ( .A1(G118), .A2(n888), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G130), .A2(n886), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(KEYINPUT114), .B(n872), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G106), .A2(n882), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G142), .A2(n883), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(n921), .ZN(n879) );
  XNOR2_X1 U979 ( .A(G162), .B(n879), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n895) );
  NAND2_X1 U981 ( .A1(G103), .A2(n882), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G139), .A2(n883), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U984 ( .A1(n886), .A2(G127), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(KEYINPUT116), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G115), .A2(n888), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n927) );
  XOR2_X1 U990 ( .A(n927), .B(G160), .Z(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U992 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n991), .B(KEYINPUT117), .ZN(n898) );
  XNOR2_X1 U994 ( .A(G171), .B(n977), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n901) );
  XOR2_X1 U996 ( .A(n899), .B(G286), .Z(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G37), .A2(n902), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n917) );
  XNOR2_X1 U1002 ( .A(G2443), .B(G2435), .ZN(n914) );
  XOR2_X1 U1003 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n906) );
  XNOR2_X1 U1004 ( .A(G2454), .B(G2430), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1006 ( .A(G2427), .B(G2438), .Z(n908) );
  XNOR2_X1 U1007 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1009 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G2451), .B(G2446), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n915), .A2(G14), .ZN(n920) );
  NAND2_X1 U1014 ( .A1(n920), .A2(G319), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n920), .ZN(G401) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n946) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G2072), .B(n927), .Z(n929) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n930), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n942) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n935), .Z(n938) );
  XOR2_X1 U1032 ( .A(G160), .B(G2084), .Z(n936) );
  XNOR2_X1 U1033 ( .A(KEYINPUT119), .B(n936), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(KEYINPUT120), .B(n943), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT52), .B(n944), .Z(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n972) );
  XNOR2_X1 U1041 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(n948), .B(KEYINPUT54), .ZN(n965) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1044 ( .A(G25), .B(n949), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(n953), .B(G27), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G2067), .B(G26), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n963), .B(KEYINPUT121), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT55), .B(n966), .ZN(n968) );
  INV_X1 U1059 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n969), .A2(G11), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT122), .B(n970), .Z(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n1027) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XOR2_X1 U1065 ( .A(G168), .B(G1966), .Z(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT57), .ZN(n995) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n977), .ZN(n983) );
  XOR2_X1 U1070 ( .A(G1956), .B(G299), .Z(n979) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G171), .B(G1961), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(n990), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1341), .B(n991), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1024) );
  INV_X1 U1084 ( .A(G16), .ZN(n1022) );
  XNOR2_X1 U1085 ( .A(n998), .B(G5), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G21), .B(G1966), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1012) );
  XOR2_X1 U1088 ( .A(G4), .B(KEYINPUT126), .Z(n1002) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1002), .B(n1001), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(KEYINPUT125), .B(G1341), .Z(n1003) );
  XNOR2_X1 U1092 ( .A(G19), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G1956), .B(G20), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1010), .Z(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G1976), .B(G23), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1025), .Z(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

