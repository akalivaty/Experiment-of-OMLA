

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586;

  XOR2_X2 U320 ( .A(n396), .B(n395), .Z(n551) );
  AND2_X1 U321 ( .A1(n571), .A2(n565), .ZN(n357) );
  NOR2_X1 U322 ( .A1(n520), .A2(n459), .ZN(n461) );
  INV_X1 U323 ( .A(KEYINPUT97), .ZN(n460) );
  XNOR2_X1 U324 ( .A(n376), .B(n345), .ZN(n350) );
  XNOR2_X1 U325 ( .A(n414), .B(n413), .ZN(n421) );
  XNOR2_X1 U326 ( .A(n444), .B(KEYINPUT126), .ZN(n584) );
  XOR2_X1 U327 ( .A(KEYINPUT64), .B(n356), .Z(n565) );
  XNOR2_X1 U328 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U329 ( .A(n388), .B(n289), .ZN(n321) );
  XOR2_X1 U330 ( .A(G169GAT), .B(KEYINPUT18), .Z(n288) );
  AND2_X1 U331 ( .A1(G226GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U332 ( .A(n429), .B(n383), .Z(n290) );
  XOR2_X1 U333 ( .A(n420), .B(n419), .Z(n291) );
  XOR2_X1 U334 ( .A(G43GAT), .B(KEYINPUT8), .Z(n292) );
  NAND2_X1 U335 ( .A1(n466), .A2(n583), .ZN(n402) );
  INV_X1 U336 ( .A(KEYINPUT21), .ZN(n314) );
  XNOR2_X1 U337 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n399) );
  OR2_X1 U338 ( .A1(n398), .A2(n397), .ZN(n400) );
  XNOR2_X1 U339 ( .A(n361), .B(G85GAT), .ZN(n345) );
  XNOR2_X1 U340 ( .A(n400), .B(n399), .ZN(n406) );
  XNOR2_X1 U341 ( .A(n317), .B(n316), .ZN(n440) );
  XNOR2_X1 U342 ( .A(n428), .B(n348), .ZN(n349) );
  INV_X1 U343 ( .A(G176GAT), .ZN(n413) );
  XNOR2_X1 U344 ( .A(n350), .B(n349), .ZN(n353) );
  XNOR2_X1 U345 ( .A(KEYINPUT26), .B(n443), .ZN(n556) );
  NOR2_X1 U346 ( .A1(n483), .A2(n556), .ZN(n444) );
  XNOR2_X1 U347 ( .A(n421), .B(n291), .ZN(n427) );
  XNOR2_X1 U348 ( .A(n401), .B(KEYINPUT36), .ZN(n466) );
  XNOR2_X1 U349 ( .A(n469), .B(KEYINPUT111), .ZN(n534) );
  INV_X1 U350 ( .A(G43GAT), .ZN(n476) );
  XNOR2_X1 U351 ( .A(n427), .B(n426), .ZN(n539) );
  XNOR2_X1 U352 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n445) );
  XNOR2_X1 U353 ( .A(n447), .B(G197GAT), .ZN(n448) );
  XNOR2_X1 U354 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n470) );
  XNOR2_X1 U355 ( .A(n476), .B(KEYINPUT40), .ZN(n477) );
  XNOR2_X1 U356 ( .A(n446), .B(n445), .ZN(G1355GAT) );
  XNOR2_X1 U357 ( .A(n449), .B(n448), .ZN(G1352GAT) );
  XNOR2_X1 U358 ( .A(n471), .B(n470), .ZN(G1336GAT) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U361 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U362 ( .A(G57GAT), .B(G1GAT), .Z(n296) );
  XNOR2_X1 U363 ( .A(G148GAT), .B(G141GAT), .ZN(n295) );
  XNOR2_X1 U364 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U365 ( .A(n298), .B(n297), .Z(n303) );
  XOR2_X1 U366 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n300) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U368 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U369 ( .A(KEYINPUT6), .B(n301), .ZN(n302) );
  XNOR2_X1 U370 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U371 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n305) );
  XNOR2_X1 U372 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n304) );
  XNOR2_X1 U373 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U374 ( .A(n307), .B(n306), .Z(n313) );
  XOR2_X1 U375 ( .A(G113GAT), .B(G127GAT), .Z(n309) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n308) );
  XNOR2_X1 U377 ( .A(n309), .B(n308), .ZN(n412) );
  XOR2_X1 U378 ( .A(G155GAT), .B(KEYINPUT3), .Z(n311) );
  XNOR2_X1 U379 ( .A(KEYINPUT88), .B(KEYINPUT2), .ZN(n310) );
  XNOR2_X1 U380 ( .A(n311), .B(n310), .ZN(n432) );
  XNOR2_X1 U381 ( .A(n412), .B(n432), .ZN(n312) );
  XOR2_X1 U382 ( .A(n313), .B(n312), .Z(n520) );
  INV_X1 U383 ( .A(KEYINPUT54), .ZN(n409) );
  XOR2_X1 U384 ( .A(G183GAT), .B(G8GAT), .Z(n364) );
  XOR2_X1 U385 ( .A(G64GAT), .B(G176GAT), .Z(n351) );
  XNOR2_X1 U386 ( .A(n364), .B(n351), .ZN(n324) );
  XNOR2_X1 U387 ( .A(G218GAT), .B(G211GAT), .ZN(n315) );
  XNOR2_X1 U388 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U389 ( .A(G197GAT), .B(G204GAT), .Z(n316) );
  XOR2_X1 U390 ( .A(KEYINPUT93), .B(n440), .Z(n320) );
  XNOR2_X1 U391 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n318) );
  XNOR2_X1 U392 ( .A(n288), .B(n318), .ZN(n422) );
  XNOR2_X1 U393 ( .A(n422), .B(G92GAT), .ZN(n319) );
  XNOR2_X1 U394 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U395 ( .A(G190GAT), .B(G36GAT), .Z(n388) );
  XOR2_X2 U396 ( .A(n324), .B(n323), .Z(n530) );
  INV_X1 U397 ( .A(n530), .ZN(n479) );
  XOR2_X1 U398 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n326) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G197GAT), .ZN(n325) );
  XNOR2_X1 U400 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .Z(n430) );
  XOR2_X1 U402 ( .A(n327), .B(n430), .Z(n330) );
  XNOR2_X1 U403 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n328) );
  XNOR2_X1 U404 ( .A(n292), .B(n328), .ZN(n383) );
  XOR2_X1 U405 ( .A(G1GAT), .B(G15GAT), .Z(n360) );
  XNOR2_X1 U406 ( .A(n383), .B(n360), .ZN(n329) );
  XNOR2_X1 U407 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n332) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U410 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U411 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U412 ( .A(G169GAT), .B(G36GAT), .Z(n336) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(G50GAT), .ZN(n335) );
  XNOR2_X1 U414 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U415 ( .A(n337), .B(KEYINPUT29), .ZN(n338) );
  XOR2_X1 U416 ( .A(n339), .B(n338), .Z(n541) );
  INV_X1 U417 ( .A(n541), .ZN(n571) );
  XOR2_X1 U418 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n341) );
  NAND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U420 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U421 ( .A(KEYINPUT31), .B(n342), .ZN(n355) );
  XOR2_X1 U422 ( .A(KEYINPUT73), .B(G99GAT), .Z(n344) );
  XNOR2_X1 U423 ( .A(KEYINPUT72), .B(G92GAT), .ZN(n343) );
  XNOR2_X1 U424 ( .A(n344), .B(n343), .ZN(n376) );
  XOR2_X1 U425 ( .A(G57GAT), .B(KEYINPUT13), .Z(n361) );
  XOR2_X1 U426 ( .A(KEYINPUT71), .B(G78GAT), .Z(n347) );
  XNOR2_X1 U427 ( .A(G148GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U428 ( .A(n347), .B(n346), .ZN(n428) );
  XOR2_X1 U429 ( .A(KEYINPUT74), .B(G204GAT), .Z(n348) );
  XOR2_X1 U430 ( .A(G120GAT), .B(G71GAT), .Z(n423) );
  XNOR2_X1 U431 ( .A(n423), .B(n351), .ZN(n352) );
  XNOR2_X1 U432 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U433 ( .A(n355), .B(n354), .Z(n580) );
  XNOR2_X1 U434 ( .A(n580), .B(KEYINPUT41), .ZN(n356) );
  XNOR2_X1 U435 ( .A(n357), .B(KEYINPUT46), .ZN(n398) );
  XOR2_X1 U436 ( .A(G211GAT), .B(G71GAT), .Z(n359) );
  XNOR2_X1 U437 ( .A(G127GAT), .B(G155GAT), .ZN(n358) );
  XNOR2_X1 U438 ( .A(n359), .B(n358), .ZN(n375) );
  XOR2_X1 U439 ( .A(n361), .B(n360), .Z(n363) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U441 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U442 ( .A(n365), .B(n364), .Z(n373) );
  XOR2_X1 U443 ( .A(KEYINPUT12), .B(G64GAT), .Z(n367) );
  XNOR2_X1 U444 ( .A(G78GAT), .B(G22GAT), .ZN(n366) );
  XNOR2_X1 U445 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U446 ( .A(KEYINPUT83), .B(KEYINPUT14), .Z(n369) );
  XNOR2_X1 U447 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n368) );
  XNOR2_X1 U448 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U449 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U450 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U451 ( .A(n375), .B(n374), .Z(n547) );
  INV_X1 U452 ( .A(n547), .ZN(n583) );
  XOR2_X1 U453 ( .A(n376), .B(G85GAT), .Z(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n378) );
  XNOR2_X1 U455 ( .A(KEYINPUT10), .B(KEYINPUT80), .ZN(n377) );
  XNOR2_X1 U456 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U457 ( .A(G106GAT), .B(KEYINPUT78), .Z(n380) );
  XNOR2_X1 U458 ( .A(G134GAT), .B(KEYINPUT67), .ZN(n379) );
  XNOR2_X1 U459 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U460 ( .A(n382), .B(n381), .Z(n394) );
  XOR2_X1 U461 ( .A(G162GAT), .B(G50GAT), .Z(n429) );
  NAND2_X1 U462 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U463 ( .A(n290), .B(n384), .ZN(n392) );
  XOR2_X1 U464 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n386) );
  XNOR2_X1 U465 ( .A(KEYINPUT81), .B(KEYINPUT79), .ZN(n385) );
  XNOR2_X1 U466 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U467 ( .A(n387), .B(KEYINPUT76), .Z(n390) );
  XNOR2_X1 U468 ( .A(n388), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U469 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U470 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U471 ( .A(n394), .B(n393), .ZN(n395) );
  INV_X1 U472 ( .A(n551), .ZN(n576) );
  OR2_X1 U473 ( .A1(n583), .A2(n576), .ZN(n397) );
  XOR2_X1 U474 ( .A(n576), .B(KEYINPUT103), .Z(n401) );
  XOR2_X1 U475 ( .A(KEYINPUT45), .B(n402), .Z(n403) );
  INV_X1 U476 ( .A(n580), .ZN(n472) );
  NAND2_X1 U477 ( .A1(n403), .A2(n472), .ZN(n404) );
  NOR2_X1 U478 ( .A1(n571), .A2(n404), .ZN(n405) );
  NOR2_X1 U479 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U480 ( .A(n407), .B(KEYINPUT48), .ZN(n555) );
  NOR2_X1 U481 ( .A1(n479), .A2(n555), .ZN(n408) );
  XNOR2_X1 U482 ( .A(n409), .B(n408), .ZN(n410) );
  NOR2_X1 U483 ( .A1(n520), .A2(n410), .ZN(n411) );
  XNOR2_X1 U484 ( .A(n411), .B(KEYINPUT65), .ZN(n483) );
  XNOR2_X1 U485 ( .A(n412), .B(G15GAT), .ZN(n414) );
  XOR2_X1 U486 ( .A(G183GAT), .B(G190GAT), .Z(n416) );
  XNOR2_X1 U487 ( .A(G99GAT), .B(G43GAT), .ZN(n415) );
  XNOR2_X1 U488 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n418) );
  XNOR2_X1 U490 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n417) );
  XNOR2_X1 U491 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U492 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U495 ( .A(n539), .ZN(n487) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n436) );
  XOR2_X1 U498 ( .A(n432), .B(KEYINPUT23), .Z(n434) );
  NAND2_X1 U499 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U501 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U502 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n438) );
  XNOR2_X1 U503 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n437) );
  XNOR2_X1 U504 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U505 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n484) );
  NAND2_X1 U507 ( .A1(n487), .A2(n484), .ZN(n443) );
  NAND2_X1 U508 ( .A1(n584), .A2(n466), .ZN(n446) );
  NAND2_X1 U509 ( .A1(n571), .A2(n584), .ZN(n449) );
  XOR2_X1 U510 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n447) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n479), .Z(n455) );
  AND2_X1 U512 ( .A1(n520), .A2(n455), .ZN(n557) );
  XNOR2_X1 U513 ( .A(n484), .B(KEYINPUT28), .ZN(n535) );
  INV_X1 U514 ( .A(n535), .ZN(n514) );
  NAND2_X1 U515 ( .A1(n557), .A2(n514), .ZN(n538) );
  XNOR2_X1 U516 ( .A(KEYINPUT94), .B(n538), .ZN(n450) );
  NOR2_X1 U517 ( .A1(n539), .A2(n450), .ZN(n451) );
  XOR2_X1 U518 ( .A(KEYINPUT95), .B(n451), .Z(n463) );
  NOR2_X1 U519 ( .A1(n487), .A2(n479), .ZN(n452) );
  NOR2_X1 U520 ( .A1(n484), .A2(n452), .ZN(n453) );
  XNOR2_X1 U521 ( .A(n453), .B(KEYINPUT25), .ZN(n457) );
  INV_X1 U522 ( .A(n556), .ZN(n454) );
  NAND2_X1 U523 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U524 ( .A1(n457), .A2(n456), .ZN(n458) );
  XOR2_X1 U525 ( .A(KEYINPUT96), .B(n458), .Z(n459) );
  XNOR2_X1 U526 ( .A(n461), .B(n460), .ZN(n462) );
  NOR2_X1 U527 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n464), .B(KEYINPUT98), .ZN(n496) );
  NOR2_X1 U529 ( .A1(n583), .A2(n496), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n465), .B(KEYINPUT104), .ZN(n467) );
  NAND2_X1 U531 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U532 ( .A(KEYINPUT37), .B(n468), .ZN(n474) );
  INV_X1 U533 ( .A(n565), .ZN(n543) );
  NOR2_X1 U534 ( .A1(n571), .A2(n543), .ZN(n517) );
  NAND2_X1 U535 ( .A1(n474), .A2(n517), .ZN(n469) );
  NAND2_X1 U536 ( .A1(n520), .A2(n534), .ZN(n471) );
  NAND2_X1 U537 ( .A1(n472), .A2(n571), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n473), .B(KEYINPUT75), .ZN(n497) );
  NAND2_X1 U539 ( .A1(n497), .A2(n474), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n475), .B(KEYINPUT38), .ZN(n513) );
  NOR2_X1 U541 ( .A1(n487), .A2(n513), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  NOR2_X1 U543 ( .A1(n479), .A2(n513), .ZN(n482) );
  INV_X1 U544 ( .A(G36GAT), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n480), .B(KEYINPUT106), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(G1329GAT) );
  NOR2_X1 U547 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(KEYINPUT55), .ZN(n486) );
  NOR2_X2 U549 ( .A1(n487), .A2(n486), .ZN(n577) );
  NAND2_X1 U550 ( .A1(n577), .A2(n565), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n491) );
  XOR2_X1 U554 ( .A(G176GAT), .B(KEYINPUT122), .Z(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1349GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n500) );
  NAND2_X1 U558 ( .A1(n551), .A2(n583), .ZN(n494) );
  XNOR2_X1 U559 ( .A(KEYINPUT16), .B(n494), .ZN(n495) );
  NOR2_X1 U560 ( .A1(n496), .A2(n495), .ZN(n518) );
  NAND2_X1 U561 ( .A1(n518), .A2(n497), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT99), .ZN(n506) );
  NAND2_X1 U563 ( .A1(n506), .A2(n520), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U565 ( .A(G1GAT), .B(n501), .Z(G1324GAT) );
  XOR2_X1 U566 ( .A(G8GAT), .B(KEYINPUT101), .Z(n503) );
  NAND2_X1 U567 ( .A1(n506), .A2(n530), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U570 ( .A1(n506), .A2(n539), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U572 ( .A1(n535), .A2(n506), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(KEYINPUT102), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(n508), .ZN(G1327GAT) );
  INV_X1 U575 ( .A(n520), .ZN(n509) );
  NOR2_X1 U576 ( .A1(n513), .A2(n509), .ZN(n512) );
  XOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  XNOR2_X1 U578 ( .A(KEYINPUT105), .B(n510), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  XNOR2_X1 U580 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n516) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1331GAT) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(n519), .Z(n526) );
  NAND2_X1 U586 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n530), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U590 ( .A(G71GAT), .B(KEYINPUT109), .Z(n525) );
  NAND2_X1 U591 ( .A1(n526), .A2(n539), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U594 ( .A1(n526), .A2(n535), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G78GAT), .B(n529), .ZN(G1335GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n534), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U599 ( .A(G99GAT), .B(KEYINPUT113), .Z(n533) );
  NAND2_X1 U600 ( .A1(n534), .A2(n539), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1338GAT) );
  NAND2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G106GAT), .ZN(G1339GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n555), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n541), .A2(n550), .ZN(n542) );
  XOR2_X1 U608 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  NOR2_X1 U609 ( .A1(n543), .A2(n550), .ZN(n545) );
  XNOR2_X1 U610 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  NOR2_X1 U613 ( .A1(n547), .A2(n550), .ZN(n548) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(n548), .Z(n549) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n554), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT117), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n569), .A2(n571), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT118), .ZN(n561) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n561), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n563) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT119), .B(n564), .Z(n567) );
  NAND2_X1 U630 ( .A1(n569), .A2(n565), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n583), .A2(n569), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U636 ( .A(G169GAT), .B(KEYINPUT121), .Z(n573) );
  NAND2_X1 U637 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(G183GAT), .B(KEYINPUT125), .Z(n575) );
  NAND2_X1 U640 ( .A1(n577), .A2(n583), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1350GAT) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1354GAT) );
endmodule

