

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U558 ( .A(KEYINPUT102), .ZN(n783) );
  XNOR2_X1 U559 ( .A(n732), .B(KEYINPUT31), .ZN(n733) );
  XNOR2_X1 U560 ( .A(n734), .B(n733), .ZN(n747) );
  NAND2_X2 U561 ( .A1(n786), .A2(n687), .ZN(n736) );
  NOR2_X1 U562 ( .A1(G651), .A2(n648), .ZN(n643) );
  NOR2_X1 U563 ( .A1(n529), .A2(n528), .ZN(n530) );
  INV_X1 U564 ( .A(G2104), .ZN(n531) );
  NOR2_X1 U565 ( .A1(G2105), .A2(n531), .ZN(n902) );
  NAND2_X1 U566 ( .A1(n902), .A2(G102), .ZN(n524) );
  XNOR2_X1 U567 ( .A(KEYINPUT85), .B(n524), .ZN(n529) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X1 U569 ( .A(KEYINPUT64), .B(n525), .Z(n526) );
  XNOR2_X2 U570 ( .A(KEYINPUT17), .B(n526), .ZN(n903) );
  NAND2_X1 U571 ( .A1(G138), .A2(n903), .ZN(n527) );
  XOR2_X1 U572 ( .A(KEYINPUT86), .B(n527), .Z(n528) );
  XNOR2_X1 U573 ( .A(n530), .B(KEYINPUT87), .ZN(n536) );
  INV_X1 U574 ( .A(G2105), .ZN(n532) );
  NOR2_X1 U575 ( .A1(n532), .A2(n531), .ZN(n906) );
  NAND2_X1 U576 ( .A1(G114), .A2(n906), .ZN(n534) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n532), .ZN(n907) );
  NAND2_X1 U578 ( .A1(G126), .A2(n907), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U580 ( .A1(n536), .A2(n535), .ZN(G164) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n634) );
  NAND2_X1 U582 ( .A1(G85), .A2(n634), .ZN(n538) );
  XOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  INV_X1 U584 ( .A(G651), .ZN(n539) );
  NOR2_X1 U585 ( .A1(n648), .A2(n539), .ZN(n632) );
  NAND2_X1 U586 ( .A1(G72), .A2(n632), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U588 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n540), .Z(n647) );
  NAND2_X1 U590 ( .A1(G60), .A2(n647), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G47), .A2(n643), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U593 ( .A1(n544), .A2(n543), .ZN(G290) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U595 ( .A1(n906), .A2(G111), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G135), .A2(n903), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n907), .A2(G123), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n902), .A2(G99), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n939) );
  XNOR2_X1 U603 ( .A(G2096), .B(n939), .ZN(n552) );
  OR2_X1 U604 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  NAND2_X1 U608 ( .A1(G89), .A2(n634), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT4), .B(n553), .Z(n554) );
  XNOR2_X1 U610 ( .A(n554), .B(KEYINPUT69), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G76), .A2(n632), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U613 ( .A(KEYINPUT5), .B(n557), .ZN(n563) );
  NAND2_X1 U614 ( .A1(G63), .A2(n647), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G51), .A2(n643), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n561) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(KEYINPUT70), .Z(n560) );
  XNOR2_X1 U618 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U620 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U623 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n837) );
  NAND2_X1 U625 ( .A1(n837), .A2(G567), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U627 ( .A1(G81), .A2(n634), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT66), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G68), .A2(n632), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(n571), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G56), .A2(n647), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n572), .Z(n575) );
  NAND2_X1 U635 ( .A1(G43), .A2(n643), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT67), .B(n573), .ZN(n574) );
  NOR2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n1003) );
  INV_X1 U639 ( .A(n1003), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n578), .A2(G860), .ZN(G153) );
  NAND2_X1 U641 ( .A1(G90), .A2(n634), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G77), .A2(n632), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT9), .B(n581), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G64), .A2(n647), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G52), .A2(n643), .ZN(n582) );
  AND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G92), .A2(n634), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G79), .A2(n632), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G66), .A2(n647), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G54), .A2(n643), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(KEYINPUT68), .B(n593), .ZN(n710) );
  INV_X1 U658 ( .A(n710), .ZN(n990) );
  NOR2_X1 U659 ( .A1(n990), .A2(G868), .ZN(n595) );
  INV_X1 U660 ( .A(G868), .ZN(n659) );
  NOR2_X1 U661 ( .A1(n659), .A2(G301), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G91), .A2(n634), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G65), .A2(n647), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G78), .A2(n632), .ZN(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT65), .B(n598), .ZN(n599) );
  NOR2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n643), .A2(G53), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(G299) );
  XNOR2_X1 U671 ( .A(KEYINPUT71), .B(G868), .ZN(n603) );
  NOR2_X1 U672 ( .A1(G286), .A2(n603), .ZN(n605) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U675 ( .A(KEYINPUT72), .B(n606), .ZN(G297) );
  INV_X1 U676 ( .A(G559), .ZN(n607) );
  NOR2_X1 U677 ( .A1(G860), .A2(n607), .ZN(n608) );
  XNOR2_X1 U678 ( .A(KEYINPUT73), .B(n608), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n609), .A2(n710), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n610), .B(KEYINPUT16), .ZN(n611) );
  XNOR2_X1 U681 ( .A(KEYINPUT74), .B(n611), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n1003), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n710), .A2(G868), .ZN(n612) );
  NOR2_X1 U684 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U685 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U686 ( .A1(G559), .A2(n710), .ZN(n657) );
  XNOR2_X1 U687 ( .A(n1003), .B(n657), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n615), .A2(G860), .ZN(n624) );
  NAND2_X1 U689 ( .A1(G67), .A2(n647), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G55), .A2(n643), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U692 ( .A(KEYINPUT76), .B(n618), .Z(n620) );
  NAND2_X1 U693 ( .A1(n632), .A2(G80), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G93), .A2(n634), .ZN(n621) );
  XNOR2_X1 U696 ( .A(KEYINPUT75), .B(n621), .ZN(n622) );
  OR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n660) );
  XOR2_X1 U698 ( .A(n624), .B(n660), .Z(G145) );
  NAND2_X1 U699 ( .A1(G62), .A2(n647), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G50), .A2(n643), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G88), .A2(n634), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G75), .A2(n632), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT79), .ZN(G303) );
  INV_X1 U707 ( .A(G303), .ZN(G166) );
  NAND2_X1 U708 ( .A1(G73), .A2(n632), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U710 ( .A1(n634), .A2(G86), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT78), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G48), .A2(n643), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G61), .A2(n647), .ZN(n638) );
  XNOR2_X1 U715 ( .A(KEYINPUT77), .B(n638), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G49), .A2(n643), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(G288) );
  XNOR2_X1 U724 ( .A(G166), .B(G305), .ZN(n653) );
  XOR2_X1 U725 ( .A(KEYINPUT19), .B(n1003), .Z(n651) );
  XNOR2_X1 U726 ( .A(G288), .B(n651), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(G299), .ZN(n656) );
  XOR2_X1 U730 ( .A(n660), .B(n656), .Z(n920) );
  XNOR2_X1 U731 ( .A(n657), .B(n920), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n666), .A2(G2072), .ZN(n667) );
  XNOR2_X1 U740 ( .A(KEYINPUT80), .B(n667), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U742 ( .A1(G69), .A2(G120), .ZN(n668) );
  NOR2_X1 U743 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U744 ( .A1(G108), .A2(n669), .ZN(n842) );
  NAND2_X1 U745 ( .A1(G567), .A2(n842), .ZN(n670) );
  XOR2_X1 U746 ( .A(KEYINPUT81), .B(n670), .Z(n675) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U749 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G96), .A2(n673), .ZN(n843) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n843), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n675), .A2(n674), .ZN(n861) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n676) );
  XNOR2_X1 U754 ( .A(KEYINPUT82), .B(n676), .ZN(n677) );
  NOR2_X1 U755 ( .A1(n861), .A2(n677), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT83), .B(n678), .Z(n841) );
  NAND2_X1 U757 ( .A1(G36), .A2(n841), .ZN(n679) );
  XNOR2_X1 U758 ( .A(n679), .B(KEYINPUT84), .ZN(G176) );
  NAND2_X1 U759 ( .A1(n906), .A2(G113), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G101), .A2(n902), .ZN(n680) );
  XOR2_X1 U761 ( .A(KEYINPUT23), .B(n680), .Z(n681) );
  NAND2_X1 U762 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U763 ( .A1(n907), .A2(G125), .ZN(n684) );
  NAND2_X1 U764 ( .A1(G137), .A2(n903), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U766 ( .A1(n686), .A2(n685), .ZN(G160) );
  INV_X1 U767 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U768 ( .A(KEYINPUT32), .B(KEYINPUT101), .ZN(n745) );
  NOR2_X2 U769 ( .A1(G164), .A2(G1384), .ZN(n786) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n785) );
  INV_X1 U771 ( .A(n785), .ZN(n687) );
  XNOR2_X1 U772 ( .A(G2078), .B(KEYINPUT25), .ZN(n962) );
  NOR2_X1 U773 ( .A1(n736), .A2(n962), .ZN(n689) );
  INV_X1 U774 ( .A(n736), .ZN(n702) );
  INV_X1 U775 ( .A(G1961), .ZN(n1009) );
  NOR2_X1 U776 ( .A1(n702), .A2(n1009), .ZN(n688) );
  NOR2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n729), .A2(G171), .ZN(n723) );
  INV_X1 U779 ( .A(KEYINPUT29), .ZN(n721) );
  INV_X1 U780 ( .A(G2072), .ZN(n932) );
  NOR2_X1 U781 ( .A1(n736), .A2(n932), .ZN(n691) );
  XNOR2_X1 U782 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n690) );
  XNOR2_X1 U783 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n736), .A2(G1956), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U786 ( .A1(G299), .A2(n695), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT28), .ZN(n719) );
  NOR2_X1 U788 ( .A1(G299), .A2(n695), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT99), .ZN(n717) );
  INV_X1 U790 ( .A(G1996), .ZN(n963) );
  NOR2_X1 U791 ( .A1(n736), .A2(n963), .ZN(n698) );
  INV_X1 U792 ( .A(KEYINPUT26), .ZN(n697) );
  XNOR2_X1 U793 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n736), .A2(G1341), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U796 ( .A1(n1003), .A2(n701), .ZN(n711) );
  OR2_X1 U797 ( .A1(n710), .A2(n711), .ZN(n715) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n702), .ZN(n703) );
  XNOR2_X1 U799 ( .A(KEYINPUT98), .B(n703), .ZN(n704) );
  NAND2_X1 U800 ( .A1(n736), .A2(G1348), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n704), .A2(n706), .ZN(n705) );
  NOR2_X1 U802 ( .A1(KEYINPUT97), .A2(n705), .ZN(n709) );
  NAND2_X1 U803 ( .A1(KEYINPUT98), .A2(KEYINPUT97), .ZN(n707) );
  NOR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U811 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n746) );
  NAND2_X1 U813 ( .A1(G8), .A2(n736), .ZN(n780) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n780), .ZN(n750) );
  NOR2_X1 U815 ( .A1(n736), .A2(G2084), .ZN(n724) );
  XNOR2_X1 U816 ( .A(n724), .B(KEYINPUT95), .ZN(n748) );
  NAND2_X1 U817 ( .A1(G8), .A2(n748), .ZN(n725) );
  NOR2_X1 U818 ( .A1(n750), .A2(n725), .ZN(n727) );
  INV_X1 U819 ( .A(KEYINPUT30), .ZN(n726) );
  XNOR2_X1 U820 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U821 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U822 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n734) );
  INV_X1 U824 ( .A(KEYINPUT100), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n746), .A2(n747), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n735), .A2(G286), .ZN(n743) );
  INV_X1 U827 ( .A(G8), .ZN(n741) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n780), .ZN(n738) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n739), .A2(G303), .ZN(n740) );
  OR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U834 ( .A(n745), .B(n744), .ZN(n770) );
  AND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n753) );
  INV_X1 U836 ( .A(n748), .ZN(n749) );
  AND2_X1 U837 ( .A1(G8), .A2(n749), .ZN(n751) );
  OR2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n768) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n983) );
  INV_X1 U841 ( .A(n983), .ZN(n754) );
  OR2_X1 U842 ( .A1(n754), .A2(n780), .ZN(n760) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n759), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n780), .A2(n755), .ZN(n764) );
  NOR2_X1 U846 ( .A1(n760), .A2(n764), .ZN(n756) );
  AND2_X1 U847 ( .A1(n768), .A2(n756), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n770), .A2(n757), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n984) );
  OR2_X1 U851 ( .A1(n760), .A2(n984), .ZN(n762) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n761) );
  AND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n998) );
  NAND2_X1 U857 ( .A1(n767), .A2(n998), .ZN(n777) );
  AND2_X1 U858 ( .A1(n768), .A2(n780), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n775) );
  INV_X1 U860 ( .A(n780), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U862 ( .A1(G8), .A2(n771), .ZN(n772) );
  OR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n782) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U867 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(n783), .ZN(n822) );
  XNOR2_X1 U871 ( .A(G1986), .B(G290), .ZN(n996) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n832) );
  NAND2_X1 U873 ( .A1(n996), .A2(n832), .ZN(n820) );
  NAND2_X1 U874 ( .A1(n902), .A2(G104), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G140), .A2(n903), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G116), .A2(n906), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G128), .A2(n907), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U883 ( .A(KEYINPUT36), .B(n795), .ZN(n891) );
  XNOR2_X1 U884 ( .A(KEYINPUT37), .B(G2067), .ZN(n830) );
  NOR2_X1 U885 ( .A1(n891), .A2(n830), .ZN(n950) );
  NAND2_X1 U886 ( .A1(n832), .A2(n950), .ZN(n828) );
  INV_X1 U887 ( .A(n828), .ZN(n818) );
  NAND2_X1 U888 ( .A1(G117), .A2(n906), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G129), .A2(n907), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n903), .A2(G141), .ZN(n798) );
  XOR2_X1 U892 ( .A(KEYINPUT90), .B(n798), .Z(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(KEYINPUT89), .Z(n802) );
  NAND2_X1 U895 ( .A1(G105), .A2(n902), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n802), .B(n801), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT91), .B(n805), .Z(n893) );
  NAND2_X1 U899 ( .A1(G1996), .A2(n893), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(KEYINPUT92), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n906), .A2(G107), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G131), .A2(n903), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U904 ( .A1(G95), .A2(n902), .ZN(n810) );
  NAND2_X1 U905 ( .A1(G119), .A2(n907), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U908 ( .A(KEYINPUT88), .B(n813), .Z(n913) );
  NAND2_X1 U909 ( .A1(n913), .A2(G1991), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n946) );
  XOR2_X1 U911 ( .A(n832), .B(KEYINPUT93), .Z(n816) );
  NAND2_X1 U912 ( .A1(n946), .A2(n816), .ZN(n817) );
  XOR2_X1 U913 ( .A(KEYINPUT94), .B(n817), .Z(n825) );
  NOR2_X1 U914 ( .A1(n818), .A2(n825), .ZN(n819) );
  AND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n835) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n893), .ZN(n937) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n913), .ZN(n942) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n942), .A2(n823), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n937), .A2(n826), .ZN(n827) );
  XNOR2_X1 U923 ( .A(KEYINPUT39), .B(n827), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n891), .A2(n830), .ZN(n943) );
  NAND2_X1 U926 ( .A1(n831), .A2(n943), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n836), .ZN(G329) );
  NAND2_X1 U930 ( .A1(n837), .A2(G2106), .ZN(n838) );
  XNOR2_X1 U931 ( .A(n838), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U933 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2090), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2084), .B(G2078), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1976), .B(G1971), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1961), .B(G1956), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(KEYINPUT41), .B(G1981), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1966), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(G229) );
  XNOR2_X1 U961 ( .A(KEYINPUT109), .B(n861), .ZN(G319) );
  XOR2_X1 U962 ( .A(G2438), .B(KEYINPUT105), .Z(n863) );
  XNOR2_X1 U963 ( .A(G1348), .B(G1341), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n873) );
  XOR2_X1 U965 ( .A(KEYINPUT106), .B(KEYINPUT103), .Z(n865) );
  XNOR2_X1 U966 ( .A(G2427), .B(G2451), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U968 ( .A(G2430), .B(KEYINPUT104), .Z(n867) );
  XNOR2_X1 U969 ( .A(G2454), .B(G2435), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U972 ( .A(G2443), .B(G2446), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n874), .A2(G14), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(KEYINPUT107), .ZN(G401) );
  NAND2_X1 U977 ( .A1(G124), .A2(n907), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n906), .A2(G112), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n902), .A2(G100), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G136), .A2(n903), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(G162) );
  NAND2_X1 U985 ( .A1(G118), .A2(n906), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G130), .A2(n907), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n902), .A2(G106), .ZN(n886) );
  NAND2_X1 U989 ( .A1(G142), .A2(n903), .ZN(n885) );
  NAND2_X1 U990 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U991 ( .A(KEYINPUT45), .B(n887), .Z(n888) );
  XNOR2_X1 U992 ( .A(KEYINPUT110), .B(n888), .ZN(n889) );
  NOR2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n896) );
  XNOR2_X1 U997 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n895) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n939), .B(n897), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(G160), .B(G162), .ZN(n898) );
  XNOR2_X1 U1001 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1002 ( .A(n901), .B(n900), .Z(n915) );
  NAND2_X1 U1003 ( .A1(n902), .A2(G103), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(G139), .A2(n903), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n906), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(G127), .A2(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT47), .B(n910), .Z(n911) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n931) );
  XNOR2_X1 U1011 ( .A(n913), .B(n931), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n916), .B(G164), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n917), .ZN(G395) );
  XOR2_X1 U1015 ( .A(KEYINPUT113), .B(G286), .Z(n919) );
  XNOR2_X1 U1016 ( .A(G171), .B(n990), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n922), .ZN(G397) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n923) );
  XOR2_X1 U1021 ( .A(KEYINPUT115), .B(n923), .Z(n924) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n924), .ZN(n928) );
  INV_X1 U1023 ( .A(G319), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n925), .A2(G401), .ZN(n926) );
  XOR2_X1 U1025 ( .A(KEYINPUT114), .B(n926), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n934) );
  XNOR2_X1 U1032 ( .A(n932), .B(n931), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1034 ( .A(KEYINPUT50), .B(n935), .Z(n953) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n938), .Z(n948) );
  XNOR2_X1 U1038 ( .A(G160), .B(G2084), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT116), .B(n951), .Z(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n954), .ZN(n956) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G29), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT117), .B(n958), .Z(n1040) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G2072), .B(G33), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n970) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n961) );
  NAND2_X1 U1056 ( .A1(n961), .A2(G28), .ZN(n968) );
  XOR2_X1 U1057 ( .A(n962), .B(G27), .Z(n965) );
  XOR2_X1 U1058 ( .A(n963), .B(G32), .Z(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT119), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n971), .ZN(n975) );
  XOR2_X1 U1064 ( .A(G34), .B(KEYINPUT120), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G2084), .B(KEYINPUT54), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(KEYINPUT118), .B(G2090), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G35), .B(n976), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT55), .B(n979), .ZN(n981) );
  INV_X1 U1072 ( .A(G29), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n982), .A2(G11), .ZN(n1038) );
  XNOR2_X1 U1075 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  NAND2_X1 U1076 ( .A1(G303), .A2(G1971), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G299), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n989), .B(KEYINPUT121), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G301), .B(G1961), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n990), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(n997), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G168), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(n1000), .B(KEYINPUT57), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G1341), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1036) );
  INV_X1 U1096 ( .A(G16), .ZN(n1034) );
  XNOR2_X1 U1097 ( .A(G5), .B(n1009), .ZN(n1028) );
  XOR2_X1 U1098 ( .A(G1956), .B(G20), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G19), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G6), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT124), .B(n1014), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(n1018), .B(KEYINPUT60), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(n1019), .B(KEYINPUT125), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(G1971), .B(G22), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(G23), .B(G1976), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(G1986), .B(G24), .Z(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(KEYINPUT58), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(G21), .B(G1966), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(KEYINPUT126), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1125 ( .A(n1041), .B(KEYINPUT127), .ZN(n1042) );
  XNOR2_X1 U1126 ( .A(KEYINPUT62), .B(n1042), .ZN(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

