

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738;

  NOR2_X1 U366 ( .A1(n613), .A2(n709), .ZN(n616) );
  NOR2_X1 U367 ( .A1(n701), .A2(n709), .ZN(n367) );
  OR2_X1 U368 ( .A1(n713), .A2(n725), .ZN(n648) );
  AND2_X1 U369 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U370 ( .A(n526), .B(KEYINPUT22), .ZN(n529) );
  INV_X1 U371 ( .A(n607), .ZN(n654) );
  AND2_X1 U372 ( .A1(n397), .A2(n347), .ZN(n396) );
  XNOR2_X1 U373 ( .A(n364), .B(KEYINPUT97), .ZN(n365) );
  AND2_X2 U374 ( .A1(n399), .A2(n402), .ZN(n348) );
  NAND2_X1 U375 ( .A1(n349), .A2(n579), .ZN(n389) );
  INV_X1 U376 ( .A(n716), .ZN(n384) );
  XNOR2_X2 U377 ( .A(n474), .B(n441), .ZN(n716) );
  NAND2_X1 U378 ( .A1(n637), .A2(n639), .ZN(n589) );
  NOR2_X1 U379 ( .A1(n621), .A2(n709), .ZN(n623) );
  NOR2_X2 U380 ( .A1(n556), .A2(n555), .ZN(n380) );
  XNOR2_X2 U381 ( .A(n389), .B(KEYINPUT39), .ZN(n611) );
  XNOR2_X2 U382 ( .A(n465), .B(G134), .ZN(n503) );
  XNOR2_X2 U383 ( .A(n399), .B(n351), .ZN(n607) );
  XNOR2_X1 U384 ( .A(n406), .B(G953), .ZN(n726) );
  XNOR2_X1 U385 ( .A(n434), .B(G113), .ZN(n435) );
  AND2_X1 U386 ( .A1(n408), .A2(n407), .ZN(n410) );
  XNOR2_X1 U387 ( .A(n387), .B(n432), .ZN(n386) );
  NAND2_X1 U388 ( .A1(n388), .A2(n605), .ZN(n387) );
  NAND2_X1 U389 ( .A1(n554), .A2(n651), .ZN(n624) );
  NOR2_X1 U390 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U391 ( .A(KEYINPUT106), .B(n531), .Z(n532) );
  NAND2_X1 U392 ( .A1(n530), .A2(n401), .ZN(n400) );
  OR2_X1 U393 ( .A1(n530), .A2(KEYINPUT67), .ZN(n404) );
  BUF_X1 U394 ( .A(n530), .Z(n651) );
  XNOR2_X1 U395 ( .A(n461), .B(n346), .ZN(n530) );
  XNOR2_X1 U396 ( .A(n506), .B(n366), .ZN(n545) );
  XNOR2_X1 U397 ( .A(n450), .B(n449), .ZN(n390) );
  XNOR2_X1 U398 ( .A(n435), .B(n436), .ZN(n438) );
  XNOR2_X1 U399 ( .A(G131), .B(KEYINPUT4), .ZN(n466) );
  XNOR2_X1 U400 ( .A(G146), .B(G125), .ZN(n343) );
  XNOR2_X2 U401 ( .A(n478), .B(n467), .ZN(n723) );
  XNOR2_X1 U402 ( .A(n516), .B(n511), .ZN(n379) );
  XNOR2_X2 U403 ( .A(n381), .B(KEYINPUT19), .ZN(n581) );
  NOR2_X2 U404 ( .A1(n609), .A2(n669), .ZN(n381) );
  NAND2_X1 U405 ( .A1(n344), .A2(n400), .ZN(n655) );
  NOR2_X1 U406 ( .A1(n571), .A2(n568), .ZN(n597) );
  OR2_X2 U407 ( .A1(n691), .A2(G902), .ZN(n430) );
  AND2_X1 U408 ( .A1(n652), .A2(KEYINPUT67), .ZN(n401) );
  XNOR2_X1 U409 ( .A(n479), .B(n423), .ZN(n661) );
  INV_X1 U410 ( .A(G472), .ZN(n423) );
  NOR2_X1 U411 ( .A1(G902), .A2(n618), .ZN(n479) );
  INV_X1 U412 ( .A(KEYINPUT8), .ZN(n449) );
  NAND2_X1 U413 ( .A1(n403), .A2(n419), .ZN(n402) );
  INV_X1 U414 ( .A(n652), .ZN(n403) );
  XNOR2_X1 U415 ( .A(G137), .B(G146), .ZN(n475) );
  INV_X1 U416 ( .A(KEYINPUT5), .ZN(n429) );
  XOR2_X1 U417 ( .A(G137), .B(G140), .Z(n467) );
  XNOR2_X1 U418 ( .A(n368), .B(n444), .ZN(n446) );
  NOR2_X1 U419 ( .A1(n385), .A2(G902), .ZN(n461) );
  XNOR2_X1 U420 ( .A(n455), .B(n359), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n454), .B(n345), .ZN(n359) );
  XNOR2_X1 U422 ( .A(G128), .B(G110), .ZN(n453) );
  XNOR2_X1 U423 ( .A(n724), .B(n467), .ZN(n457) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n569) );
  INV_X1 U425 ( .A(KEYINPUT28), .ZN(n356) );
  INV_X1 U426 ( .A(KEYINPUT75), .ZN(n573) );
  XNOR2_X1 U427 ( .A(G478), .B(KEYINPUT102), .ZN(n366) );
  NAND2_X1 U428 ( .A1(n505), .A2(n504), .ZN(n506) );
  INV_X1 U429 ( .A(G902), .ZN(n504) );
  INV_X1 U430 ( .A(n661), .ZN(n542) );
  BUF_X1 U431 ( .A(n726), .Z(n372) );
  XNOR2_X1 U432 ( .A(n413), .B(n417), .ZN(n702) );
  XNOR2_X1 U433 ( .A(n415), .B(n414), .ZN(n413) );
  XNOR2_X1 U434 ( .A(n500), .B(n502), .ZN(n414) );
  AND2_X2 U435 ( .A1(n375), .A2(n392), .ZN(n705) );
  INV_X1 U436 ( .A(n648), .ZN(n371) );
  NOR2_X1 U437 ( .A1(n372), .A2(G952), .ZN(n709) );
  NOR2_X1 U438 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U439 ( .A1(KEYINPUT47), .A2(n668), .ZN(n590) );
  INV_X1 U440 ( .A(KEYINPUT17), .ZN(n369) );
  OR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n484) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n534) );
  INV_X1 U443 ( .A(KEYINPUT66), .ZN(n373) );
  XOR2_X1 U444 ( .A(KEYINPUT69), .B(G119), .Z(n452) );
  NOR2_X1 U445 ( .A1(n725), .A2(n354), .ZN(n407) );
  XNOR2_X1 U446 ( .A(G146), .B(G101), .ZN(n468) );
  XNOR2_X1 U447 ( .A(G107), .B(G104), .ZN(n439) );
  NAND2_X1 U448 ( .A1(G237), .A2(G234), .ZN(n489) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n612) );
  XNOR2_X1 U450 ( .A(n464), .B(n463), .ZN(n652) );
  XNOR2_X1 U451 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n517) );
  XNOR2_X1 U452 ( .A(n474), .B(n427), .ZN(n477) );
  XNOR2_X1 U453 ( .A(n476), .B(n428), .ZN(n427) );
  XNOR2_X1 U454 ( .A(n475), .B(n429), .ZN(n428) );
  INV_X1 U455 ( .A(KEYINPUT64), .ZN(n406) );
  XNOR2_X1 U456 ( .A(n472), .B(n370), .ZN(n441) );
  XNOR2_X1 U457 ( .A(n440), .B(G122), .ZN(n370) );
  INV_X1 U458 ( .A(KEYINPUT16), .ZN(n440) );
  XNOR2_X1 U459 ( .A(n503), .B(n416), .ZN(n415) );
  XNOR2_X1 U460 ( .A(n501), .B(n499), .ZN(n416) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(G140), .Z(n510) );
  XNOR2_X1 U462 ( .A(G104), .B(G131), .ZN(n509) );
  XNOR2_X1 U463 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U464 ( .A(G143), .B(G122), .ZN(n513) );
  XNOR2_X1 U465 ( .A(n481), .B(n480), .ZN(n684) );
  AND2_X1 U466 ( .A1(n537), .A2(n600), .ZN(n481) );
  NOR2_X1 U467 ( .A1(n684), .A2(n541), .ZN(n498) );
  INV_X1 U468 ( .A(n651), .ZN(n567) );
  INV_X1 U469 ( .A(KEYINPUT107), .ZN(n422) );
  NAND2_X1 U470 ( .A1(n394), .A2(n400), .ZN(n393) );
  XNOR2_X1 U471 ( .A(n538), .B(KEYINPUT89), .ZN(n541) );
  INV_X1 U472 ( .A(n600), .ZN(n382) );
  XNOR2_X1 U473 ( .A(n363), .B(n420), .ZN(n385) );
  XNOR2_X1 U474 ( .A(n421), .B(n451), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n457), .B(n358), .ZN(n363) );
  XNOR2_X1 U476 ( .A(n391), .B(n352), .ZN(n613) );
  NAND2_X1 U477 ( .A1(n705), .A2(G210), .ZN(n391) );
  INV_X1 U478 ( .A(KEYINPUT40), .ZN(n361) );
  INV_X1 U479 ( .A(n592), .ZN(n424) );
  INV_X1 U480 ( .A(KEYINPUT119), .ZN(n377) );
  XNOR2_X1 U481 ( .A(n698), .B(n697), .ZN(n699) );
  AND2_X1 U482 ( .A1(n404), .A2(n402), .ZN(n344) );
  XOR2_X1 U483 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n345) );
  XOR2_X1 U484 ( .A(n460), .B(n459), .Z(n346) );
  OR2_X1 U485 ( .A1(n400), .A2(KEYINPUT95), .ZN(n347) );
  AND2_X1 U486 ( .A1(n418), .A2(n578), .ZN(n349) );
  AND2_X1 U487 ( .A1(n402), .A2(KEYINPUT95), .ZN(n350) );
  INV_X1 U488 ( .A(KEYINPUT67), .ZN(n419) );
  XOR2_X1 U489 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n351) );
  XOR2_X1 U490 ( .A(n448), .B(n447), .Z(n352) );
  XNOR2_X1 U491 ( .A(n723), .B(n431), .ZN(n691) );
  OR2_X1 U492 ( .A1(n647), .A2(n612), .ZN(n353) );
  AND2_X1 U493 ( .A1(n612), .A2(n412), .ZN(n354) );
  OR2_X1 U494 ( .A1(n612), .A2(n412), .ZN(n355) );
  NAND2_X1 U495 ( .A1(n597), .A2(n575), .ZN(n357) );
  NOR2_X2 U496 ( .A1(n552), .A2(n532), .ZN(n533) );
  XNOR2_X2 U497 ( .A(n533), .B(KEYINPUT32), .ZN(n737) );
  NOR2_X2 U498 ( .A1(n735), .A2(n738), .ZN(n580) );
  XNOR2_X2 U499 ( .A(n362), .B(n361), .ZN(n735) );
  XNOR2_X2 U500 ( .A(n559), .B(n558), .ZN(n713) );
  NAND2_X1 U501 ( .A1(n371), .A2(KEYINPUT2), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n360), .B(KEYINPUT83), .ZN(n554) );
  NAND2_X1 U503 ( .A1(n553), .A2(n654), .ZN(n360) );
  NAND2_X1 U504 ( .A1(n409), .A2(n353), .ZN(n375) );
  XNOR2_X1 U505 ( .A(n445), .B(n369), .ZN(n368) );
  NAND2_X1 U506 ( .A1(n611), .A2(n635), .ZN(n362) );
  NAND2_X1 U507 ( .A1(n507), .A2(n508), .ZN(n364) );
  NOR2_X2 U508 ( .A1(n698), .A2(G902), .ZN(n518) );
  XNOR2_X2 U509 ( .A(n544), .B(G475), .ZN(n523) );
  XNOR2_X2 U510 ( .A(n518), .B(n517), .ZN(n544) );
  XNOR2_X2 U511 ( .A(n365), .B(n379), .ZN(n698) );
  XNOR2_X1 U512 ( .A(n367), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U513 ( .A(n702), .ZN(n505) );
  OR2_X2 U514 ( .A1(n724), .A2(KEYINPUT11), .ZN(n507) );
  NOR2_X2 U515 ( .A1(n737), .A2(n630), .ZN(n535) );
  NOR2_X2 U516 ( .A1(n655), .A2(n654), .ZN(n537) );
  XNOR2_X2 U517 ( .A(n430), .B(G469), .ZN(n399) );
  NAND2_X1 U518 ( .A1(n736), .A2(n522), .ZN(n374) );
  XNOR2_X2 U519 ( .A(n456), .B(KEYINPUT10), .ZN(n724) );
  XNOR2_X1 U520 ( .A(n376), .B(KEYINPUT105), .ZN(n525) );
  NAND2_X1 U521 ( .A1(n671), .A2(n652), .ZN(n376) );
  XNOR2_X1 U522 ( .A(n378), .B(n377), .ZN(G63) );
  NOR2_X2 U523 ( .A1(n704), .A2(n709), .ZN(n378) );
  NOR2_X2 U524 ( .A1(n546), .A2(n545), .ZN(n635) );
  NAND2_X1 U525 ( .A1(n380), .A2(n557), .ZN(n559) );
  NAND2_X2 U526 ( .A1(n383), .A2(n382), .ZN(n552) );
  INV_X1 U527 ( .A(n529), .ZN(n383) );
  NAND2_X1 U528 ( .A1(n483), .A2(n612), .ZN(n488) );
  XNOR2_X2 U529 ( .A(n384), .B(n446), .ZN(n483) );
  XNOR2_X1 U530 ( .A(n385), .B(n707), .ZN(n708) );
  NAND2_X1 U531 ( .A1(n386), .A2(n433), .ZN(n725) );
  XNOR2_X1 U532 ( .A(n580), .B(KEYINPUT46), .ZN(n388) );
  XNOR2_X1 U533 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U534 ( .A1(n390), .A2(G221), .ZN(n421) );
  NAND2_X1 U535 ( .A1(n390), .A2(G217), .ZN(n417) );
  NAND2_X1 U536 ( .A1(n396), .A2(n393), .ZN(n572) );
  AND2_X1 U537 ( .A1(n395), .A2(n404), .ZN(n394) );
  AND2_X1 U538 ( .A1(n399), .A2(n350), .ZN(n395) );
  NAND2_X1 U539 ( .A1(n398), .A2(n405), .ZN(n397) );
  NAND2_X1 U540 ( .A1(n348), .A2(n404), .ZN(n398) );
  INV_X1 U541 ( .A(KEYINPUT95), .ZN(n405) );
  OR2_X1 U542 ( .A1(n713), .A2(n355), .ZN(n411) );
  NAND2_X1 U543 ( .A1(n713), .A2(n412), .ZN(n408) );
  NAND2_X1 U544 ( .A1(n410), .A2(n411), .ZN(n409) );
  INV_X1 U545 ( .A(KEYINPUT79), .ZN(n412) );
  NAND2_X1 U546 ( .A1(n579), .A2(n578), .ZN(n585) );
  INV_X1 U547 ( .A(n673), .ZN(n418) );
  XNOR2_X1 U548 ( .A(n661), .B(n422), .ZN(n575) );
  NAND2_X1 U549 ( .A1(n424), .A2(n589), .ZN(n583) );
  NAND2_X1 U550 ( .A1(n424), .A2(n631), .ZN(n632) );
  NAND2_X1 U551 ( .A1(n424), .A2(n635), .ZN(n636) );
  NAND2_X1 U552 ( .A1(n426), .A2(n425), .ZN(n592) );
  INV_X1 U553 ( .A(n581), .ZN(n425) );
  INV_X1 U554 ( .A(n582), .ZN(n426) );
  XNOR2_X2 U555 ( .A(n438), .B(n437), .ZN(n474) );
  XNOR2_X2 U556 ( .A(n503), .B(n466), .ZN(n478) );
  XNOR2_X2 U557 ( .A(G143), .B(G128), .ZN(n465) );
  XNOR2_X1 U558 ( .A(n472), .B(n471), .ZN(n431) );
  XNOR2_X1 U559 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X2 U560 ( .A1(n523), .A2(n545), .ZN(n524) );
  XNOR2_X2 U561 ( .A(G146), .B(G125), .ZN(n456) );
  XNOR2_X1 U562 ( .A(KEYINPUT48), .B(KEYINPUT81), .ZN(n432) );
  AND2_X1 U563 ( .A1(n646), .A2(n644), .ZN(n433) );
  XNOR2_X1 U564 ( .A(n465), .B(KEYINPUT18), .ZN(n443) );
  INV_X2 U565 ( .A(KEYINPUT3), .ZN(n434) );
  XNOR2_X1 U566 ( .A(n470), .B(n469), .ZN(n471) );
  INV_X1 U567 ( .A(KEYINPUT23), .ZN(n451) );
  INV_X1 U568 ( .A(KEYINPUT82), .ZN(n551) );
  XNOR2_X1 U569 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U570 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U571 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U572 ( .A(KEYINPUT116), .B(KEYINPUT54), .Z(n448) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(G119), .ZN(n436) );
  XNOR2_X1 U574 ( .A(G116), .B(G101), .ZN(n437) );
  XNOR2_X1 U575 ( .A(n439), .B(G110), .ZN(n472) );
  NAND2_X1 U576 ( .A1(G224), .A2(n726), .ZN(n442) );
  XNOR2_X1 U577 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U578 ( .A(n343), .B(KEYINPUT4), .Z(n445) );
  XNOR2_X1 U579 ( .A(n483), .B(KEYINPUT55), .ZN(n447) );
  NAND2_X1 U580 ( .A1(n726), .A2(G234), .ZN(n450) );
  XNOR2_X1 U581 ( .A(n452), .B(n453), .ZN(n455) );
  XOR2_X1 U582 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n454) );
  XOR2_X1 U583 ( .A(KEYINPUT76), .B(KEYINPUT25), .Z(n460) );
  NAND2_X1 U584 ( .A1(n612), .A2(G234), .ZN(n458) );
  XNOR2_X1 U585 ( .A(n458), .B(KEYINPUT20), .ZN(n462) );
  NAND2_X1 U586 ( .A1(n462), .A2(G217), .ZN(n459) );
  XOR2_X1 U587 ( .A(KEYINPUT21), .B(KEYINPUT94), .Z(n464) );
  NAND2_X1 U588 ( .A1(G221), .A2(n462), .ZN(n463) );
  NAND2_X1 U589 ( .A1(n726), .A2(G227), .ZN(n470) );
  XNOR2_X1 U590 ( .A(n468), .B(KEYINPUT90), .ZN(n469) );
  NOR2_X2 U591 ( .A1(G237), .A2(G953), .ZN(n473) );
  XNOR2_X1 U592 ( .A(n473), .B(KEYINPUT74), .ZN(n512) );
  NAND2_X1 U593 ( .A1(n512), .A2(G210), .ZN(n476) );
  XNOR2_X1 U594 ( .A(n478), .B(n477), .ZN(n618) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(n542), .ZN(n600) );
  XNOR2_X1 U596 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n480) );
  NAND2_X1 U597 ( .A1(G214), .A2(n484), .ZN(n482) );
  XOR2_X1 U598 ( .A(KEYINPUT86), .B(n482), .Z(n669) );
  XOR2_X1 U599 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n486) );
  NAND2_X1 U600 ( .A1(G210), .A2(n484), .ZN(n485) );
  XNOR2_X1 U601 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X2 U602 ( .A(n488), .B(n487), .ZN(n609) );
  INV_X1 U603 ( .A(G953), .ZN(n649) );
  XNOR2_X1 U604 ( .A(n489), .B(KEYINPUT14), .ZN(n490) );
  NAND2_X1 U605 ( .A1(G952), .A2(n490), .ZN(n682) );
  NOR2_X1 U606 ( .A1(G953), .A2(n682), .ZN(n564) );
  INV_X1 U607 ( .A(n564), .ZN(n494) );
  NAND2_X1 U608 ( .A1(n490), .A2(G902), .ZN(n491) );
  XOR2_X1 U609 ( .A(KEYINPUT87), .B(n491), .Z(n561) );
  INV_X1 U610 ( .A(n561), .ZN(n492) );
  NOR2_X1 U611 ( .A1(G898), .A2(n649), .ZN(n718) );
  NAND2_X1 U612 ( .A1(n492), .A2(n718), .ZN(n493) );
  NAND2_X1 U613 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U614 ( .A(KEYINPUT88), .B(n495), .Z(n496) );
  NOR2_X2 U615 ( .A1(n581), .A2(n496), .ZN(n497) );
  XNOR2_X2 U616 ( .A(n497), .B(KEYINPUT0), .ZN(n538) );
  XNOR2_X1 U617 ( .A(n498), .B(KEYINPUT34), .ZN(n520) );
  XOR2_X1 U618 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n500) );
  XNOR2_X1 U619 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n499) );
  XOR2_X1 U620 ( .A(G122), .B(KEYINPUT99), .Z(n502) );
  XNOR2_X1 U621 ( .A(G107), .B(G116), .ZN(n501) );
  NAND2_X1 U622 ( .A1(n724), .A2(KEYINPUT11), .ZN(n508) );
  XOR2_X1 U623 ( .A(n510), .B(n509), .Z(n511) );
  NAND2_X1 U624 ( .A1(G214), .A2(n512), .ZN(n515) );
  XNOR2_X1 U625 ( .A(n513), .B(G113), .ZN(n514) );
  NAND2_X1 U626 ( .A1(n545), .A2(n523), .ZN(n584) );
  XNOR2_X1 U627 ( .A(n584), .B(KEYINPUT77), .ZN(n519) );
  XNOR2_X2 U628 ( .A(n521), .B(KEYINPUT35), .ZN(n736) );
  INV_X1 U629 ( .A(KEYINPUT44), .ZN(n522) );
  XNOR2_X2 U630 ( .A(n524), .B(KEYINPUT104), .ZN(n671) );
  NAND2_X1 U631 ( .A1(n525), .A2(n538), .ZN(n526) );
  NOR2_X1 U632 ( .A1(n575), .A2(n529), .ZN(n527) );
  NAND2_X1 U633 ( .A1(n527), .A2(n567), .ZN(n528) );
  NOR2_X1 U634 ( .A1(n607), .A2(n528), .ZN(n630) );
  NOR2_X1 U635 ( .A1(n654), .A2(n651), .ZN(n531) );
  NAND2_X1 U636 ( .A1(n534), .A2(n535), .ZN(n557) );
  NAND2_X1 U637 ( .A1(n535), .A2(n736), .ZN(n536) );
  NAND2_X1 U638 ( .A1(n536), .A2(KEYINPUT44), .ZN(n550) );
  XOR2_X1 U639 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n540) );
  AND2_X1 U640 ( .A1(n537), .A2(n661), .ZN(n664) );
  NAND2_X1 U641 ( .A1(n664), .A2(n538), .ZN(n539) );
  XNOR2_X1 U642 ( .A(n540), .B(n539), .ZN(n640) );
  NOR2_X1 U643 ( .A1(n541), .A2(n572), .ZN(n543) );
  NAND2_X1 U644 ( .A1(n543), .A2(n542), .ZN(n626) );
  NAND2_X1 U645 ( .A1(n640), .A2(n626), .ZN(n547) );
  XOR2_X1 U646 ( .A(G475), .B(n544), .Z(n546) );
  INV_X1 U647 ( .A(n635), .ZN(n637) );
  NAND2_X1 U648 ( .A1(n546), .A2(n545), .ZN(n639) );
  NAND2_X1 U649 ( .A1(n547), .A2(n589), .ZN(n548) );
  XOR2_X1 U650 ( .A(n548), .B(KEYINPUT103), .Z(n549) );
  NAND2_X1 U651 ( .A1(n550), .A2(n549), .ZN(n556) );
  INV_X1 U652 ( .A(n624), .ZN(n555) );
  INV_X1 U653 ( .A(KEYINPUT45), .ZN(n558) );
  INV_X1 U654 ( .A(n609), .ZN(n586) );
  XNOR2_X1 U655 ( .A(KEYINPUT38), .B(n586), .ZN(n673) );
  INV_X1 U656 ( .A(n669), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n576), .A2(n671), .ZN(n667) );
  NOR2_X1 U658 ( .A1(n673), .A2(n667), .ZN(n560) );
  XNOR2_X1 U659 ( .A(KEYINPUT41), .B(n560), .ZN(n683) );
  NOR2_X1 U660 ( .A1(n372), .A2(n561), .ZN(n562) );
  XOR2_X1 U661 ( .A(KEYINPUT108), .B(n562), .Z(n563) );
  NOR2_X1 U662 ( .A1(G900), .A2(n563), .ZN(n565) );
  NOR2_X1 U663 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U664 ( .A(KEYINPUT78), .B(n566), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n652), .A2(n567), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n569), .A2(n399), .ZN(n582) );
  NOR2_X1 U667 ( .A1(n683), .A2(n582), .ZN(n570) );
  XNOR2_X1 U668 ( .A(n570), .B(KEYINPUT42), .ZN(n738) );
  AND2_X1 U669 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U670 ( .A(KEYINPUT30), .B(n577), .ZN(n578) );
  NAND2_X1 U671 ( .A1(n583), .A2(KEYINPUT47), .ZN(n588) );
  NOR2_X1 U672 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n634) );
  NAND2_X1 U674 ( .A1(n588), .A2(n634), .ZN(n595) );
  INV_X1 U675 ( .A(n589), .ZN(n668) );
  XNOR2_X1 U676 ( .A(n590), .B(KEYINPUT73), .ZN(n591) );
  XNOR2_X1 U677 ( .A(n593), .B(KEYINPUT72), .ZN(n594) );
  NOR2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U679 ( .A(KEYINPUT71), .B(n596), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n597), .A2(n635), .ZN(n598) );
  NOR2_X1 U681 ( .A1(n669), .A2(n598), .ZN(n599) );
  NAND2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n609), .A2(n606), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n601), .B(KEYINPUT36), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n602), .A2(n607), .ZN(n643) );
  INV_X1 U686 ( .A(n643), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  OR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U689 ( .A(KEYINPUT43), .B(n608), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n646) );
  INV_X1 U691 ( .A(n639), .ZN(n631) );
  NAND2_X1 U692 ( .A1(n631), .A2(n611), .ZN(n644) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n647) );
  XOR2_X1 U694 ( .A(KEYINPUT80), .B(KEYINPUT117), .Z(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(KEYINPUT56), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n616), .B(n615), .ZN(G51) );
  NAND2_X1 U697 ( .A1(n705), .A2(G472), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT62), .B(KEYINPUT109), .Z(n617) );
  XOR2_X1 U699 ( .A(KEYINPUT63), .B(KEYINPUT110), .Z(n622) );
  XNOR2_X1 U700 ( .A(n623), .B(n622), .ZN(G57) );
  XNOR2_X1 U701 ( .A(G101), .B(n624), .ZN(G3) );
  NOR2_X1 U702 ( .A1(n637), .A2(n626), .ZN(n625) );
  XOR2_X1 U703 ( .A(G104), .B(n625), .Z(G6) );
  NOR2_X1 U704 ( .A1(n639), .A2(n626), .ZN(n628) );
  XNOR2_X1 U705 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U707 ( .A(G107), .B(n629), .ZN(G9) );
  XOR2_X1 U708 ( .A(G110), .B(n630), .Z(G12) );
  XOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .Z(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(G30) );
  XNOR2_X1 U711 ( .A(G143), .B(n634), .ZN(G45) );
  XNOR2_X1 U712 ( .A(n636), .B(G146), .ZN(G48) );
  NOR2_X1 U713 ( .A1(n640), .A2(n637), .ZN(n638) );
  XOR2_X1 U714 ( .A(G113), .B(n638), .Z(G15) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U716 ( .A(G116), .B(n641), .Z(G18) );
  XOR2_X1 U717 ( .A(G125), .B(KEYINPUT37), .Z(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G134), .B(n644), .ZN(G36) );
  XOR2_X1 U720 ( .A(G140), .B(KEYINPUT111), .Z(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(G42) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n689) );
  NOR2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT49), .B(n653), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT50), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT112), .B(n657), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U731 ( .A(KEYINPUT113), .B(n662), .Z(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(KEYINPUT51), .B(n665), .Z(n666) );
  NOR2_X1 U734 ( .A1(n683), .A2(n666), .ZN(n678) );
  INV_X1 U735 ( .A(n667), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n684), .A2(n676), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U742 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U743 ( .A(KEYINPUT52), .B(n680), .ZN(n681) );
  NOR2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U747 ( .A(n687), .B(KEYINPUT115), .ZN(n688) );
  NOR2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U749 ( .A(KEYINPUT53), .B(n690), .ZN(G75) );
  XNOR2_X1 U750 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n691), .B(KEYINPUT57), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U753 ( .A1(n705), .A2(G469), .ZN(n694) );
  XOR2_X1 U754 ( .A(n695), .B(n694), .Z(n696) );
  NOR2_X1 U755 ( .A1(n709), .A2(n696), .ZN(G54) );
  NAND2_X1 U756 ( .A1(n705), .A2(G475), .ZN(n700) );
  INV_X1 U757 ( .A(KEYINPUT59), .ZN(n697) );
  NAND2_X1 U758 ( .A1(G478), .A2(n705), .ZN(n703) );
  XNOR2_X1 U759 ( .A(n702), .B(n703), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n705), .A2(G217), .ZN(n706) );
  XNOR2_X1 U761 ( .A(n706), .B(KEYINPUT120), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n710) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n711), .A2(G898), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT121), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n713), .A2(G953), .ZN(n714) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n722) );
  XNOR2_X1 U769 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT122), .B(n716), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n722), .B(n721), .ZN(G69) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n728) );
  XNOR2_X1 U775 ( .A(n728), .B(n725), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(n372), .ZN(n732) );
  XNOR2_X1 U777 ( .A(G227), .B(n728), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U781 ( .A(KEYINPUT125), .B(n733), .Z(G72) );
  XOR2_X1 U782 ( .A(G131), .B(KEYINPUT126), .Z(n734) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(G33) );
  XNOR2_X1 U784 ( .A(G122), .B(n736), .ZN(G24) );
  XOR2_X1 U785 ( .A(n737), .B(G119), .Z(G21) );
  XOR2_X1 U786 ( .A(G137), .B(n738), .Z(G39) );
endmodule

