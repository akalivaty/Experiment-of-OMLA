//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G97), .A2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G77), .A2(G244), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n207), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n216), .B2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G13), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n221), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n218), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G226), .B(G232), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n251), .A4(new_n252), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT73), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT73), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n253), .B2(new_n254), .ZN(new_n259));
  OAI21_X1  g0059(.A(G107), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT75), .ZN(new_n261));
  XOR2_X1   g0061(.A(G97), .B(G107), .Z(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT6), .A2(G97), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n262), .A2(KEYINPUT6), .B1(G107), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT75), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(G107), .C1(new_n257), .C2(new_n259), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G77), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n261), .A2(new_n265), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G97), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n271), .A2(new_n226), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n279), .B(new_n275), .C1(G1), .C2(new_n249), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n278), .B1(new_n280), .B2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G244), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT4), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n284), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G283), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT67), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n227), .A2(new_n295), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT5), .A2(G41), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT5), .A2(G41), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n304), .A2(G257), .A3(new_n293), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n298), .A2(new_n299), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n306), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n310), .B(new_n307), .C1(new_n291), .C2(new_n297), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(G200), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n273), .A2(new_n282), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n298), .A2(new_n314), .A3(new_n306), .A4(new_n308), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n311), .B2(G169), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n273), .B2(new_n282), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  OAI211_X1 g0120(.A(G226), .B(new_n284), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(G232), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n297), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n293), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G238), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n297), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n328), .A2(new_n305), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n327), .A2(new_n330), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n325), .B2(new_n326), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n330), .A4(new_n331), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G169), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(G179), .A3(new_n339), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(new_n345), .A3(G169), .A4(new_n341), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G68), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G20), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n251), .A2(G33), .ZN(new_n350));
  INV_X1    g0150(.A(G77), .ZN(new_n351));
  INV_X1    g0151(.A(new_n268), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n349), .B1(new_n350), .B2(new_n351), .C1(new_n352), .C2(new_n202), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n272), .B1(new_n274), .B2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n275), .A2(G68), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT11), .B1(new_n353), .B2(new_n272), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n347), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT8), .B(G58), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n276), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n356), .B2(new_n366), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(G226), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n370));
  OAI211_X1 g0170(.A(G223), .B(new_n284), .C1(new_n319), .C2(new_n320), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G87), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n370), .A2(new_n371), .A3(new_n375), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n297), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n332), .B1(new_n329), .B2(G232), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(G190), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n257), .B2(new_n259), .ZN(new_n380));
  INV_X1    g0180(.A(G58), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n348), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n201), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n268), .A2(G159), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n319), .A2(new_n320), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n388), .B2(new_n251), .ZN(new_n389));
  INV_X1    g0189(.A(new_n256), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n272), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n369), .B(new_n379), .C1(new_n387), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n377), .A2(new_n378), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT17), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n258), .B1(new_n389), .B2(new_n390), .ZN(new_n400));
  INV_X1    g0200(.A(new_n259), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n348), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n385), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n392), .A2(new_n272), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n368), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n396), .A4(new_n379), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n377), .A2(G179), .A3(new_n378), .ZN(new_n410));
  INV_X1    g0210(.A(G169), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n377), .B2(new_n378), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n405), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n369), .B1(new_n387), .B2(new_n393), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(KEYINPUT18), .C1(new_n412), .C2(new_n410), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n275), .A2(G77), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n356), .A2(new_n351), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n366), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n421));
  XOR2_X1   g0221(.A(KEYINPUT15), .B(G87), .Z(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n350), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n419), .B(new_n420), .C1(new_n424), .C2(new_n272), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n426));
  INV_X1    g0226(.A(G107), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n283), .A2(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G238), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n426), .B1(new_n427), .B2(new_n283), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n297), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n329), .A2(G244), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n333), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT68), .B1(new_n433), .B2(G179), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n332), .B1(new_n430), .B2(new_n297), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT68), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n314), .A4(new_n432), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n425), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n411), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n364), .A2(new_n418), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT9), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n203), .A2(G20), .ZN(new_n444));
  INV_X1    g0244(.A(G150), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n444), .B1(new_n445), .B2(new_n352), .C1(new_n350), .C2(new_n365), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n272), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n276), .A2(new_n202), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n355), .A2(G50), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT69), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(KEYINPUT69), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n443), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n453), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n451), .A3(KEYINPUT9), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n458));
  INV_X1    g0258(.A(G223), .ZN(new_n459));
  OAI221_X1 g0259(.A(new_n458), .B1(new_n351), .B2(new_n283), .C1(new_n428), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n297), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n329), .A2(G226), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n333), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G190), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT70), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n463), .B2(G200), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n457), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT10), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT10), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n457), .A2(new_n470), .A3(new_n465), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n450), .B1(new_n463), .B2(G179), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n411), .B2(new_n463), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n433), .A2(G200), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n425), .C1(new_n299), .C2(new_n433), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n340), .A2(G200), .A3(new_n341), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n335), .A2(G190), .A3(new_n339), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n361), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n442), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n304), .A2(G264), .A3(new_n293), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(new_n284), .C1(new_n319), .C2(new_n320), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT80), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n283), .A2(new_n486), .A3(G250), .A4(new_n284), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G294), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n485), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n483), .B1(new_n490), .B2(new_n297), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n299), .A3(new_n306), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT81), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n306), .ZN(new_n494));
  INV_X1    g0294(.A(G200), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(new_n497), .A3(new_n299), .A4(new_n306), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G116), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G20), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n251), .A2(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT23), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(new_n250), .B2(new_n252), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G87), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n251), .B(G87), .C1(new_n319), .C2(new_n320), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n502), .B(new_n504), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT24), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n283), .A2(new_n505), .A3(new_n251), .A4(G87), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n501), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n504), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n279), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT25), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n275), .B2(G107), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n275), .A2(new_n518), .A3(G107), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n280), .A2(new_n427), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n499), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n490), .A2(new_n297), .ZN(new_n525));
  INV_X1    g0325(.A(new_n483), .ZN(new_n526));
  AND4_X1   g0326(.A1(G179), .A2(new_n525), .A3(new_n306), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n411), .B1(new_n491), .B2(new_n306), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n517), .B2(new_n522), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n514), .A2(new_n515), .A3(new_n504), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n515), .B1(new_n514), .B2(new_n504), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n272), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n522), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(KEYINPUT79), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n529), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n275), .A2(G116), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n280), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n290), .B(new_n251), .C1(G33), .C2(new_n277), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT78), .ZN(new_n543));
  AOI221_X4 g0343(.A(new_n543), .B1(new_n540), .B2(G20), .C1(new_n271), .C2(new_n226), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT78), .B1(new_n272), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(KEYINPUT20), .B(new_n542), .C1(new_n544), .C2(new_n546), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n539), .B(new_n541), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n283), .A2(G257), .A3(new_n284), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n283), .A2(G264), .A3(G1698), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n388), .A2(G303), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n297), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n304), .A2(new_n293), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G270), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n558), .A3(new_n306), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G169), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n538), .B1(new_n551), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n549), .A2(new_n550), .ZN(new_n562));
  INV_X1    g0362(.A(new_n539), .ZN(new_n563));
  INV_X1    g0363(.A(new_n541), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n555), .A2(new_n297), .B1(new_n557), .B2(G270), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n411), .B1(new_n566), .B2(new_n306), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(KEYINPUT21), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n559), .A2(new_n314), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n561), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n559), .A2(G200), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n566), .A2(G190), .A3(new_n306), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n551), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G244), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n575));
  OAI211_X1 g0375(.A(G238), .B(new_n284), .C1(new_n319), .C2(new_n320), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n500), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n297), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n301), .A2(G274), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n580), .A2(G250), .A3(new_n293), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n422), .A2(new_n275), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(new_n251), .A3(G33), .A4(G97), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n209), .B1(new_n323), .B2(new_n251), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n589), .B2(new_n586), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n251), .B(G68), .C1(new_n319), .C2(new_n320), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT77), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n283), .A2(new_n593), .A3(new_n251), .A4(G68), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n585), .B1(new_n595), .B2(new_n272), .ZN(new_n596));
  INV_X1    g0396(.A(new_n280), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G87), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n578), .A2(G190), .A3(new_n579), .A4(new_n582), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n584), .A2(new_n596), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n422), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n583), .A2(new_n411), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n578), .A2(new_n314), .A3(new_n579), .A4(new_n582), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n574), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n537), .A2(new_n571), .A3(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n318), .A2(new_n482), .A3(new_n524), .A4(new_n607), .ZN(G372));
  AND3_X1   g0408(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n596), .A2(KEYINPUT82), .A3(new_n598), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT82), .B1(new_n596), .B2(new_n598), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n584), .A2(new_n599), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n528), .A2(new_n527), .B1(new_n517), .B2(new_n522), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n615), .A2(new_n561), .A3(new_n568), .A4(new_n570), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n318), .A2(new_n524), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n317), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(new_n605), .ZN(new_n620));
  INV_X1    g0420(.A(new_n317), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n605), .A2(new_n600), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT26), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n482), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(KEYINPUT83), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n441), .A2(new_n481), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n363), .A2(new_n627), .B1(new_n398), .B2(new_n407), .ZN(new_n628));
  INV_X1    g0428(.A(new_n417), .ZN(new_n629));
  OR3_X1    g0429(.A1(new_n628), .A2(KEYINPUT84), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT84), .B1(new_n628), .B2(new_n629), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n472), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n475), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(new_n633), .ZN(G369));
  INV_X1    g0434(.A(new_n574), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n221), .A2(G20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n274), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT85), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT27), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n551), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n571), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n571), .A2(new_n646), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n635), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g0449(.A(KEYINPUT86), .B(G330), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n571), .A2(new_n645), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n531), .A2(new_n536), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n529), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n524), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n524), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n537), .A2(new_n644), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n659), .B2(new_n652), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n527), .ZN(new_n663));
  INV_X1    g0463(.A(new_n528), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n534), .B2(new_n535), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n645), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(G399));
  NAND4_X1  g0469(.A1(new_n607), .A2(new_n318), .A3(new_n524), .A4(new_n645), .ZN(new_n670));
  INV_X1    g0470(.A(new_n583), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n491), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT88), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n307), .B1(new_n291), .B2(new_n297), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT88), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n675), .A3(new_n491), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n569), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n676), .A2(new_n674), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n569), .A4(new_n673), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n494), .A2(new_n314), .A3(new_n559), .A4(new_n583), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(new_n311), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n644), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(KEYINPUT31), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n650), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n281), .B1(new_n270), .B2(new_n272), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(new_n622), .A3(new_n316), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n618), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n317), .A2(new_n614), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n609), .B1(new_n694), .B2(KEYINPUT26), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n318), .A2(new_n524), .A3(new_n614), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n537), .A2(new_n571), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n693), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n690), .B1(new_n698), .B2(new_n645), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n624), .A2(new_n690), .A3(new_n645), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n689), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n274), .ZN(new_n703));
  INV_X1    g0503(.A(new_n223), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT87), .B1(new_n704), .B2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n704), .A2(KEYINPUT87), .A3(G41), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G1), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n588), .A2(new_n209), .A3(new_n540), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n710), .A2(new_n711), .B1(new_n229), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n703), .A2(new_n713), .ZN(G364));
  XNOR2_X1  g0514(.A(new_n651), .B(KEYINPUT89), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n274), .B1(new_n636), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n715), .B(new_n719), .C1(new_n650), .C2(new_n649), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n251), .A2(G179), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G190), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(KEYINPUT92), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(KEYINPUT92), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n495), .A2(G190), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n727), .A2(G329), .B1(G283), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  NOR2_X1   g0532(.A1(new_n251), .A2(new_n314), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G190), .A3(new_n495), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G322), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n299), .A2(new_n495), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n721), .ZN(new_n738));
  INV_X1    g0538(.A(G303), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n388), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n733), .A2(new_n728), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G317), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT33), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(KEYINPUT33), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n733), .A2(new_n737), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G326), .ZN(new_n749));
  INV_X1    g0549(.A(G294), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n299), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n251), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n746), .B(new_n749), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n733), .A2(new_n722), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n740), .B(new_n753), .C1(G311), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n732), .A2(new_n736), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n351), .ZN(new_n758));
  INV_X1    g0558(.A(new_n738), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G87), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n760), .B(new_n283), .C1(new_n427), .C2(new_n729), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT91), .Z(new_n762));
  INV_X1    g0562(.A(new_n723), .ZN(new_n763));
  XNOR2_X1  g0563(.A(KEYINPUT90), .B(G159), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT32), .Z(new_n766));
  INV_X1    g0566(.A(new_n752), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G97), .B1(new_n748), .B2(G50), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n735), .A2(G58), .B1(new_n742), .B2(G68), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n762), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n757), .B1(new_n758), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n226), .B1(G20), .B2(new_n411), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n283), .B1(new_n243), .B2(G45), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G45), .B2(new_n229), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n283), .A2(G355), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n223), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n772), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G116), .B2(new_n704), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n771), .A2(new_n772), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n779), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n649), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n720), .B1(new_n719), .B2(new_n785), .ZN(G396));
  NOR2_X1   g0586(.A1(new_n440), .A2(new_n644), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n425), .A2(new_n642), .A3(new_n643), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n439), .A2(new_n438), .B1(new_n788), .B2(new_n477), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n624), .B2(new_n645), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n273), .A2(new_n282), .A3(new_n312), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n524), .B(new_n792), .C1(new_n691), .C2(new_n316), .ZN(new_n793));
  INV_X1    g0593(.A(new_n614), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n571), .A2(new_n665), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n619), .B(new_n605), .C1(new_n618), .C2(new_n692), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n645), .B(new_n790), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT95), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n624), .A2(KEYINPUT95), .A3(new_n645), .A4(new_n790), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n791), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(new_n689), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n719), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n772), .A2(new_n777), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G137), .A2(new_n748), .B1(new_n755), .B2(new_n764), .ZN(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n808), .B2(new_n734), .C1(new_n445), .C2(new_n741), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n388), .B1(new_n727), .B2(G132), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n730), .A2(G68), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n767), .A2(G58), .B1(new_n759), .B2(G50), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n388), .B1(new_n734), .B2(new_n750), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n747), .A2(new_n739), .B1(new_n741), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G97), .C2(new_n767), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n427), .A2(new_n738), .B1(new_n754), .B2(new_n540), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n727), .B2(G311), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(new_n209), .C2(new_n729), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n772), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n718), .B1(G77), .B2(new_n806), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT94), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n778), .B2(new_n790), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n804), .A2(new_n826), .ZN(G384));
  INV_X1    g0627(.A(KEYINPUT39), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n395), .A2(G169), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n377), .A2(G179), .A3(new_n378), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n830), .A3(new_n642), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n415), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n403), .A2(new_n404), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n833), .A2(new_n369), .A3(new_n396), .A4(new_n379), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT98), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n832), .A2(new_n834), .A3(new_n838), .A4(new_n835), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n348), .B1(new_n255), .B2(new_n256), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n399), .B1(new_n841), .B2(new_n385), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n404), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n369), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n831), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n835), .B1(new_n845), .B2(new_n834), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n642), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n418), .A2(new_n849), .A3(new_n844), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  INV_X1    g0652(.A(new_n844), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n642), .B(new_n853), .C1(new_n408), .C2(new_n417), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n846), .B1(new_n837), .B2(new_n839), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n851), .A2(new_n856), .A3(KEYINPUT99), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(new_n852), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n828), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT102), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n848), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n850), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n408), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n398), .A2(new_n407), .A3(KEYINPUT101), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n417), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n415), .A3(new_n849), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n832), .A2(new_n834), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n840), .B1(new_n835), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n852), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n860), .B1(new_n874), .B2(new_n828), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT97), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n363), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n347), .A2(KEYINPUT97), .A3(new_n362), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(new_n644), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n629), .A2(new_n642), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n644), .A2(new_n362), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n481), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n347), .A2(KEYINPUT97), .A3(new_n362), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT97), .B1(new_n347), .B2(new_n362), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n364), .A2(new_n644), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n800), .A2(new_n801), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n787), .B(KEYINPUT96), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n859), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT100), .B1(new_n857), .B2(new_n859), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n889), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n881), .A2(new_n882), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n701), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n482), .B1(new_n699), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n633), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n897), .B(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n862), .A2(new_n863), .B1(new_n872), .B2(new_n852), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n686), .A2(new_n687), .A3(new_n790), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n889), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n904), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n894), .B2(new_n895), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n908), .B2(new_n905), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n482), .A2(new_n688), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n650), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n901), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n274), .B2(new_n636), .ZN(new_n914));
  OAI211_X1 g0714(.A(G20), .B(new_n227), .C1(new_n264), .C2(KEYINPUT35), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n540), .B(new_n915), .C1(KEYINPUT35), .C2(new_n264), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT36), .Z(new_n917));
  OAI21_X1  g0717(.A(G77), .B1(new_n381), .B2(new_n348), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n918), .A2(new_n229), .B1(G50), .B2(new_n348), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G1), .A3(new_n221), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n914), .A2(new_n917), .A3(new_n920), .ZN(G367));
  XOR2_X1   g0721(.A(new_n708), .B(KEYINPUT41), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n661), .B1(new_n715), .B2(new_n660), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n924), .A2(new_n689), .A3(new_n700), .A4(new_n701), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n621), .A2(new_n792), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n691), .A2(new_n645), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n621), .A2(new_n645), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n931), .C2(new_n668), .ZN(new_n932));
  NAND2_X1  g0732(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n933));
  OR2_X1    g0733(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n930), .A2(new_n667), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT45), .B1(new_n931), .B2(new_n668), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT45), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n930), .A2(new_n938), .A3(new_n667), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n662), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n661), .A2(KEYINPUT107), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n940), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n932), .B(new_n935), .C1(new_n937), .C2(new_n939), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n941), .A3(new_n662), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n925), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n923), .B1(new_n947), .B2(new_n702), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(KEYINPUT108), .B(new_n923), .C1(new_n947), .C2(new_n702), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n716), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n645), .A2(new_n612), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n609), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n794), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT103), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n930), .B(KEYINPUT104), .ZN(new_n959));
  INV_X1    g0759(.A(new_n537), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n644), .B1(new_n961), .B2(new_n621), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n656), .A2(new_n926), .A3(new_n927), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT42), .Z(new_n964));
  OAI221_X1 g0764(.A(new_n956), .B1(KEYINPUT105), .B2(new_n958), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n959), .A2(new_n662), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n958), .A2(KEYINPUT105), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n965), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n952), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n234), .A2(new_n704), .A3(new_n283), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n781), .B(new_n971), .C1(new_n704), .C2(new_n422), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT109), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n718), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n748), .A2(G143), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n759), .A2(G58), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n742), .A2(new_n764), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n283), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n735), .A2(G150), .B1(new_n763), .B2(G137), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n202), .B2(new_n754), .C1(new_n351), .C2(new_n729), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(G68), .C2(new_n767), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n735), .A2(G303), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n729), .A2(new_n277), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G283), .B2(new_n755), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n743), .B2(new_n723), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n767), .A2(G107), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n759), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n748), .A2(G311), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT46), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n738), .B2(new_n540), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n388), .B1(new_n741), .B2(new_n750), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n985), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n981), .B1(new_n982), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n974), .B1(new_n995), .B2(new_n772), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n972), .A2(new_n973), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n955), .A2(new_n784), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n970), .A2(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n924), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n702), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(new_n925), .A3(new_n708), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G322), .A2(new_n748), .B1(new_n755), .B2(G303), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n742), .A2(G311), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n743), .C2(new_n734), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n1008));
  AOI22_X1  g0808(.A1(new_n1007), .A2(new_n1008), .B1(G283), .B2(new_n767), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n750), .B2(new_n738), .C1(new_n1008), .C2(new_n1007), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n763), .A2(G326), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n283), .B1(new_n730), .B2(G116), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n735), .A2(G50), .B1(new_n759), .B2(G77), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n348), .B2(new_n754), .ZN(new_n1018));
  XOR2_X1   g0818(.A(KEYINPUT111), .B(G150), .Z(new_n1019));
  AOI211_X1 g0819(.A(new_n983), .B(new_n1018), .C1(new_n763), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n742), .A2(new_n366), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n423), .A2(new_n752), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G159), .B2(new_n748), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n283), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n719), .B1(new_n1025), .B2(new_n772), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n239), .A2(new_n300), .A3(new_n283), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n365), .A2(G50), .ZN(new_n1028));
  XOR2_X1   g0828(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1029));
  AOI21_X1  g0829(.A(G45), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n348), .B2(new_n351), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n711), .B1(new_n1031), .B2(new_n388), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n223), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n780), .C1(new_n427), .C2(new_n223), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1026), .B(new_n1034), .C1(new_n659), .C2(new_n784), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1003), .B(new_n1035), .C1(new_n716), .C2(new_n1001), .ZN(G393));
  NOR2_X1   g0836(.A1(new_n223), .A2(new_n277), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n704), .A2(new_n283), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n781), .B(new_n1037), .C1(new_n246), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n388), .B1(new_n730), .B2(G87), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n348), .B2(new_n738), .C1(new_n808), .C2(new_n723), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1042));
  INV_X1    g0842(.A(G159), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n734), .A2(new_n1043), .B1(new_n747), .B2(new_n445), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT51), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n767), .A2(G77), .B1(new_n742), .B2(G50), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n366), .B2(new_n755), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n752), .A2(new_n540), .B1(new_n741), .B2(new_n739), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT114), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n750), .C2(new_n754), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT115), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n735), .A2(G311), .B1(new_n748), .B2(G317), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n388), .B1(new_n729), .B2(new_n427), .C1(new_n816), .C2(new_n738), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n763), .A2(G322), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n718), .B1(new_n1061), .B2(new_n823), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1039), .B(new_n1062), .C1(new_n959), .C2(new_n779), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n944), .A2(new_n946), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n717), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n944), .A2(new_n925), .A3(new_n946), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n708), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1065), .B1(new_n1067), .B2(new_n947), .ZN(G390));
  INV_X1    g0868(.A(new_n880), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n698), .A2(new_n645), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1070), .A2(new_n789), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n787), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n879), .A2(new_n884), .B1(new_n364), .B2(new_n644), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n874), .B(new_n1069), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n880), .B1(new_n893), .B2(new_n889), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n875), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n686), .A2(new_n687), .A3(G330), .A4(new_n790), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT117), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT117), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n889), .A2(new_n903), .A3(new_n1080), .A4(G330), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1077), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n891), .B1(new_n800), .B2(new_n801), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1069), .B1(new_n1084), .B2(new_n1073), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n860), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT116), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n686), .A2(new_n687), .A3(new_n650), .A4(new_n790), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1073), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1087), .B(new_n1074), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1083), .A2(new_n1091), .A3(new_n717), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n283), .B1(new_n754), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G132), .B2(new_n735), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n767), .A2(G159), .B1(new_n742), .B2(G137), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n1096), .C1(new_n1097), .C2(new_n726), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n759), .A2(new_n1019), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT53), .Z(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n747), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1098), .B(new_n1102), .C1(G50), .C2(new_n730), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G283), .A2(new_n748), .B1(new_n742), .B2(G107), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n283), .B1(new_n767), .B2(G77), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n760), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n812), .B1(new_n277), .B2(new_n754), .C1(new_n726), .C2(new_n750), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G116), .C2(new_n735), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n772), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n718), .B1(new_n366), .B2(new_n806), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT118), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n875), .C2(new_n778), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1092), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(KEYINPUT119), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(KEYINPUT119), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n482), .A2(G330), .A3(new_n688), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n899), .A2(new_n1117), .A3(new_n475), .A4(new_n632), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1073), .A2(new_n1089), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1079), .A2(new_n1081), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n893), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1090), .A2(new_n1072), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1118), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1116), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1083), .A2(new_n1091), .A3(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n708), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1114), .A2(new_n1115), .A3(new_n1128), .ZN(G378));
  INV_X1    g0929(.A(new_n1118), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n874), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n857), .A2(new_n859), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT100), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n859), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n904), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n1132), .C1(new_n1137), .C2(KEYINPUT40), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n452), .A2(new_n453), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT55), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n472), .A2(new_n1140), .A3(new_n475), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n472), .B2(new_n475), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1139), .B(new_n849), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n849), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1141), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1144), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1138), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n908), .A2(new_n905), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1156), .A2(G330), .A3(new_n1132), .A4(new_n1153), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1155), .A2(new_n897), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n897), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1131), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n881), .A2(new_n882), .A3(new_n896), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1157), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1153), .B1(new_n909), .B2(G330), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1155), .A2(new_n897), .A3(new_n1157), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(KEYINPUT57), .A3(new_n1131), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1162), .A2(new_n1169), .A3(new_n708), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1154), .A2(new_n777), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n805), .A2(new_n202), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n752), .A2(new_n445), .B1(new_n747), .B2(new_n1097), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g0974(.A(G137), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1175), .A2(new_n754), .B1(new_n738), .B2(new_n1093), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G132), .B2(new_n742), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1174), .B(new_n1177), .C1(new_n1101), .C2(new_n734), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT59), .Z(new_n1179));
  AOI21_X1  g0979(.A(G41), .B1(new_n763), .B2(G124), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G33), .B1(new_n730), .B2(new_n764), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n202), .B1(new_n319), .B2(G41), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n734), .A2(new_n427), .B1(new_n729), .B2(new_n381), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n727), .B2(G283), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n755), .A2(new_n422), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n747), .A2(new_n540), .B1(new_n741), .B2(new_n277), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G68), .B2(new_n767), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G41), .B(new_n283), .C1(new_n759), .C2(G77), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT58), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1182), .A2(new_n1183), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n719), .B1(new_n1192), .B2(new_n772), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1171), .A2(new_n1172), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1168), .B2(new_n717), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1170), .A2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n717), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n388), .B1(new_n729), .B2(new_n351), .C1(new_n277), .C2(new_n738), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1022), .B(new_n1200), .C1(G294), .C2(new_n748), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n735), .A2(G283), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n427), .A2(new_n754), .B1(new_n741), .B2(new_n540), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT122), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n727), .A2(G303), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n388), .B1(new_n730), .B2(G58), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n202), .B2(new_n752), .C1(new_n445), .C2(new_n754), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G128), .B2(new_n727), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n748), .A2(G132), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n1175), .B2(new_n734), .C1(new_n741), .C2(new_n1093), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1209), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n738), .A2(new_n1043), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1206), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1217), .A2(new_n772), .B1(new_n348), .B2(new_n805), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n718), .B(new_n1218), .C1(new_n889), .C2(new_n778), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1199), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT124), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1199), .A2(KEYINPUT124), .A3(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1121), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1125), .A2(new_n1225), .A3(new_n923), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1170), .A3(new_n1196), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT125), .Z(new_n1231));
  NOR3_X1   g1031(.A1(new_n1229), .A2(G387), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G390), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1224), .A4(new_n1226), .ZN(G407));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n643), .A2(G213), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1166), .A2(KEYINPUT126), .A3(new_n1167), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n716), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1131), .B(new_n923), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1194), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1237), .B1(new_n1244), .B2(new_n1228), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1236), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n709), .B1(new_n1225), .B2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(new_n1125), .C1(new_n1247), .C2(new_n1225), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1224), .A2(G384), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G384), .B1(new_n1224), .B2(new_n1249), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G2897), .B(new_n1237), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1252), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1237), .A2(G2897), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1250), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT61), .B1(new_n1246), .B2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1236), .A2(new_n1245), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1236), .A2(new_n1245), .A3(new_n1263), .A4(new_n1260), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1259), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G390), .B1(new_n970), .B2(new_n999), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n999), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1267), .B(new_n1233), .C1(new_n952), .C2(new_n969), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT127), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(G396), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(KEYINPUT127), .B(new_n1270), .C1(new_n1266), .C2(new_n1268), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1236), .A2(new_n1245), .A3(new_n1260), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1274), .B1(new_n1276), .B2(KEYINPUT63), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1257), .B1(new_n1236), .B2(new_n1245), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1261), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1275), .A2(new_n1282), .ZN(G405));
  NAND3_X1  g1083(.A1(new_n1274), .A2(new_n1229), .A3(new_n1236), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1236), .A2(new_n1229), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1284), .A2(new_n1286), .A3(new_n1260), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1260), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G402));
endmodule


