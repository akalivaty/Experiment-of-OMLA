

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G2104), .A2(n555), .ZN(n899) );
  OR2_X1 U554 ( .A1(n719), .A2(n1012), .ZN(n720) );
  NOR2_X1 U555 ( .A1(n721), .A2(n720), .ZN(n727) );
  NOR2_X1 U556 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U557 ( .A1(n603), .A2(n602), .ZN(n1012) );
  XOR2_X2 U558 ( .A(KEYINPUT1), .B(n576), .Z(n609) );
  INV_X1 U559 ( .A(n915), .ZN(n991) );
  XNOR2_X1 U560 ( .A(n791), .B(n790), .ZN(n801) );
  NAND2_X1 U561 ( .A1(n527), .A2(n523), .ZN(n791) );
  NAND2_X1 U562 ( .A1(n780), .A2(n779), .ZN(n792) );
  AND2_X1 U563 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U564 ( .A1(n727), .A2(n991), .ZN(n728) );
  NOR2_X1 U565 ( .A1(n560), .A2(n559), .ZN(G164) );
  BUF_X1 U566 ( .A(n637), .Z(n638) );
  NAND2_X2 U567 ( .A1(n535), .A2(n531), .ZN(n898) );
  NOR2_X1 U568 ( .A1(G543), .A2(n575), .ZN(n576) );
  NAND2_X1 U569 ( .A1(G160), .A2(G40), .ZN(n802) );
  NOR2_X1 U570 ( .A1(n772), .A2(n541), .ZN(n540) );
  XNOR2_X1 U571 ( .A(n771), .B(KEYINPUT32), .ZN(n780) );
  AND2_X1 U572 ( .A1(n549), .A2(n845), .ZN(n548) );
  OR2_X1 U573 ( .A1(n524), .A2(KEYINPUT106), .ZN(n549) );
  NAND2_X1 U574 ( .A1(n533), .A2(KEYINPUT65), .ZN(n535) );
  NAND2_X1 U575 ( .A1(n532), .A2(n534), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XNOR2_X1 U577 ( .A(n910), .B(n526), .ZN(n911) );
  XNOR2_X1 U578 ( .A(n538), .B(KEYINPUT30), .ZN(n754) );
  NAND2_X1 U579 ( .A1(n536), .A2(n537), .ZN(n539) );
  INV_X1 U580 ( .A(G1966), .ZN(n537) );
  INV_X1 U581 ( .A(G2084), .ZN(n525) );
  NOR2_X1 U582 ( .A1(G164), .A2(G1384), .ZN(n803) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  INV_X1 U584 ( .A(KEYINPUT65), .ZN(n534) );
  INV_X1 U585 ( .A(KEYINPUT33), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n786), .A2(n785), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n801), .A2(n522), .ZN(n543) );
  NAND2_X1 U588 ( .A1(n548), .A2(n520), .ZN(n545) );
  AND2_X1 U589 ( .A1(n521), .A2(n547), .ZN(n544) );
  INV_X1 U590 ( .A(KEYINPUT106), .ZN(n547) );
  XNOR2_X1 U591 ( .A(KEYINPUT68), .B(G543), .ZN(n571) );
  AND2_X2 U592 ( .A1(n555), .A2(G2104), .ZN(n902) );
  XNOR2_X1 U593 ( .A(n551), .B(n550), .ZN(n553) );
  NOR2_X1 U594 ( .A1(n568), .A2(n569), .ZN(G160) );
  NAND2_X1 U595 ( .A1(n524), .A2(KEYINPUT106), .ZN(n520) );
  NOR2_X2 U596 ( .A1(G651), .A2(n683), .ZN(n610) );
  NOR2_X2 U597 ( .A1(n575), .A2(n683), .ZN(n606) );
  AND2_X1 U598 ( .A1(n800), .A2(n799), .ZN(n521) );
  BUF_X1 U599 ( .A(n731), .Z(n763) );
  AND2_X1 U600 ( .A1(n521), .A2(n548), .ZN(n522) );
  NOR2_X1 U601 ( .A1(n789), .A2(n788), .ZN(n523) );
  NOR2_X1 U602 ( .A1(n831), .A2(n830), .ZN(n524) );
  INV_X1 U603 ( .A(G8), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G160), .B(n525), .ZN(n949) );
  INV_X1 U605 ( .A(G160), .ZN(n526) );
  NAND2_X1 U606 ( .A1(n529), .A2(n528), .ZN(n527) );
  XNOR2_X1 U607 ( .A(n530), .B(KEYINPUT64), .ZN(n529) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n538) );
  INV_X1 U609 ( .A(n798), .ZN(n536) );
  INV_X1 U610 ( .A(n539), .ZN(n776) );
  NAND2_X1 U611 ( .A1(n546), .A2(n542), .ZN(n846) );
  NAND2_X1 U612 ( .A1(n543), .A2(n545), .ZN(n542) );
  NAND2_X1 U613 ( .A1(n801), .A2(n544), .ZN(n546) );
  NOR2_X1 U614 ( .A1(G2105), .A2(G2104), .ZN(n556) );
  INV_X1 U615 ( .A(G2105), .ZN(n555) );
  NOR2_X1 U616 ( .A1(n763), .A2(n868), .ZN(n722) );
  INV_X1 U617 ( .A(KEYINPUT98), .ZN(n737) );
  XNOR2_X1 U618 ( .A(n738), .B(n737), .ZN(n741) );
  NAND2_X1 U619 ( .A1(n715), .A2(n803), .ZN(n731) );
  INV_X1 U620 ( .A(n1007), .ZN(n789) );
  INV_X1 U621 ( .A(KEYINPUT105), .ZN(n790) );
  INV_X1 U622 ( .A(KEYINPUT15), .ZN(n615) );
  INV_X1 U623 ( .A(KEYINPUT87), .ZN(n550) );
  XNOR2_X1 U624 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U625 ( .A(KEYINPUT0), .ZN(n570) );
  INV_X1 U626 ( .A(KEYINPUT23), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n571), .B(n570), .ZN(n683) );
  XNOR2_X1 U628 ( .A(n565), .B(n564), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n898), .A2(G114), .ZN(n551) );
  NAND2_X1 U630 ( .A1(n899), .A2(G126), .ZN(n552) );
  NAND2_X1 U631 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U632 ( .A(n554), .B(KEYINPUT88), .ZN(n560) );
  NAND2_X1 U633 ( .A1(G102), .A2(n902), .ZN(n558) );
  XOR2_X1 U634 ( .A(KEYINPUT17), .B(n556), .Z(n637) );
  NAND2_X1 U635 ( .A1(G138), .A2(n637), .ZN(n557) );
  NAND2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U637 ( .A1(G125), .A2(n899), .ZN(n562) );
  NAND2_X1 U638 ( .A1(G137), .A2(n637), .ZN(n561) );
  NAND2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n569) );
  NAND2_X1 U640 ( .A1(G113), .A2(n898), .ZN(n563) );
  XNOR2_X1 U641 ( .A(n563), .B(KEYINPUT66), .ZN(n567) );
  NAND2_X1 U642 ( .A1(G101), .A2(n902), .ZN(n565) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U644 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U645 ( .A1(G651), .A2(G543), .ZN(n671) );
  NAND2_X1 U646 ( .A1(G90), .A2(n671), .ZN(n573) );
  INV_X1 U647 ( .A(G651), .ZN(n575) );
  NAND2_X1 U648 ( .A1(G77), .A2(n606), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U650 ( .A(n574), .B(KEYINPUT9), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G64), .A2(n609), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U653 ( .A1(G52), .A2(n610), .ZN(n579) );
  XNOR2_X1 U654 ( .A(KEYINPUT69), .B(n579), .ZN(n580) );
  NOR2_X1 U655 ( .A1(n581), .A2(n580), .ZN(G171) );
  AND2_X1 U656 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U657 ( .A(G57), .ZN(G237) );
  NAND2_X1 U658 ( .A1(n671), .A2(G89), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U660 ( .A1(G76), .A2(n606), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT5), .ZN(n590) );
  NAND2_X1 U663 ( .A1(G63), .A2(n609), .ZN(n587) );
  NAND2_X1 U664 ( .A1(G51), .A2(n610), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U666 ( .A(KEYINPUT6), .B(n588), .Z(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n591), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U669 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U670 ( .A1(G7), .A2(G661), .ZN(n592) );
  XOR2_X1 U671 ( .A(n592), .B(KEYINPUT10), .Z(n937) );
  NAND2_X1 U672 ( .A1(n937), .A2(G567), .ZN(n593) );
  XOR2_X1 U673 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  NAND2_X1 U674 ( .A1(n671), .A2(G81), .ZN(n594) );
  XNOR2_X1 U675 ( .A(n594), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U676 ( .A1(G68), .A2(n606), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n598) );
  XOR2_X1 U678 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n597) );
  XNOR2_X1 U679 ( .A(n598), .B(n597), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n609), .A2(G56), .ZN(n599) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n599), .Z(n600) );
  NAND2_X1 U682 ( .A1(n610), .A2(G43), .ZN(n602) );
  XNOR2_X1 U683 ( .A(G860), .B(KEYINPUT71), .ZN(n629) );
  NOR2_X1 U684 ( .A1(n1012), .A2(n629), .ZN(n604) );
  XOR2_X1 U685 ( .A(KEYINPUT72), .B(n604), .Z(G153) );
  INV_X1 U686 ( .A(G868), .ZN(n686) );
  NOR2_X1 U687 ( .A1(n686), .A2(G171), .ZN(n605) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT73), .ZN(n619) );
  NAND2_X1 U689 ( .A1(G92), .A2(n671), .ZN(n608) );
  NAND2_X1 U690 ( .A1(G79), .A2(n606), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G66), .A2(n609), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G54), .A2(n610), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT74), .B(n617), .Z(n915) );
  NAND2_X1 U697 ( .A1(n686), .A2(n915), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(G284) );
  NAND2_X1 U699 ( .A1(G65), .A2(n609), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G53), .A2(n610), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G91), .A2(n671), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G78), .A2(n606), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n994) );
  INV_X1 U706 ( .A(n994), .ZN(G299) );
  NOR2_X1 U707 ( .A1(G868), .A2(G299), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT75), .B(n626), .Z(n628) );
  NOR2_X1 U709 ( .A1(G286), .A2(n686), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(G297) );
  NAND2_X1 U711 ( .A1(n629), .A2(G559), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n630), .A2(n991), .ZN(n631) );
  XNOR2_X1 U713 ( .A(n631), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U714 ( .A1(G868), .A2(n1012), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n991), .A2(G868), .ZN(n632) );
  NOR2_X1 U716 ( .A1(G559), .A2(n632), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(G282) );
  NAND2_X1 U718 ( .A1(G123), .A2(n899), .ZN(n635) );
  XNOR2_X1 U719 ( .A(n635), .B(KEYINPUT18), .ZN(n636) );
  XNOR2_X1 U720 ( .A(n636), .B(KEYINPUT76), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G135), .A2(n638), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n641), .B(KEYINPUT77), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G111), .A2(n898), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n902), .A2(G99), .ZN(n644) );
  XOR2_X1 U727 ( .A(KEYINPUT78), .B(n644), .Z(n645) );
  NOR2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n948) );
  XNOR2_X1 U729 ( .A(n948), .B(G2096), .ZN(n647) );
  INV_X1 U730 ( .A(G2100), .ZN(n865) );
  NAND2_X1 U731 ( .A1(n647), .A2(n865), .ZN(G156) );
  NAND2_X1 U732 ( .A1(G93), .A2(n671), .ZN(n649) );
  NAND2_X1 U733 ( .A1(G67), .A2(n609), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n606), .A2(G80), .ZN(n650) );
  XOR2_X1 U736 ( .A(KEYINPUT80), .B(n650), .Z(n651) );
  NOR2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n610), .A2(G55), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n691) );
  NAND2_X1 U740 ( .A1(n991), .A2(G559), .ZN(n655) );
  XNOR2_X1 U741 ( .A(n1012), .B(n655), .ZN(n694) );
  NOR2_X1 U742 ( .A1(G860), .A2(n694), .ZN(n656) );
  XOR2_X1 U743 ( .A(KEYINPUT79), .B(n656), .Z(n657) );
  XOR2_X1 U744 ( .A(n691), .B(n657), .Z(G145) );
  NAND2_X1 U745 ( .A1(G88), .A2(n671), .ZN(n659) );
  NAND2_X1 U746 ( .A1(G75), .A2(n606), .ZN(n658) );
  NAND2_X1 U747 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U748 ( .A1(G62), .A2(n609), .ZN(n661) );
  NAND2_X1 U749 ( .A1(G50), .A2(n610), .ZN(n660) );
  NAND2_X1 U750 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U751 ( .A1(n663), .A2(n662), .ZN(G166) );
  INV_X1 U752 ( .A(G166), .ZN(G303) );
  NAND2_X1 U753 ( .A1(G72), .A2(n606), .ZN(n665) );
  NAND2_X1 U754 ( .A1(G47), .A2(n610), .ZN(n664) );
  NAND2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U756 ( .A1(G85), .A2(n671), .ZN(n666) );
  XNOR2_X1 U757 ( .A(KEYINPUT67), .B(n666), .ZN(n667) );
  NOR2_X1 U758 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U759 ( .A1(n609), .A2(G60), .ZN(n669) );
  NAND2_X1 U760 ( .A1(n670), .A2(n669), .ZN(G290) );
  NAND2_X1 U761 ( .A1(G86), .A2(n671), .ZN(n673) );
  NAND2_X1 U762 ( .A1(G61), .A2(n609), .ZN(n672) );
  NAND2_X1 U763 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U764 ( .A1(n606), .A2(G73), .ZN(n674) );
  XOR2_X1 U765 ( .A(KEYINPUT2), .B(n674), .Z(n675) );
  NOR2_X1 U766 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U767 ( .A1(n610), .A2(G48), .ZN(n677) );
  NAND2_X1 U768 ( .A1(n678), .A2(n677), .ZN(G305) );
  NAND2_X1 U769 ( .A1(G49), .A2(n610), .ZN(n680) );
  NAND2_X1 U770 ( .A1(G74), .A2(G651), .ZN(n679) );
  NAND2_X1 U771 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U772 ( .A1(n609), .A2(n681), .ZN(n682) );
  XOR2_X1 U773 ( .A(KEYINPUT81), .B(n682), .Z(n685) );
  NAND2_X1 U774 ( .A1(G87), .A2(n683), .ZN(n684) );
  NAND2_X1 U775 ( .A1(n685), .A2(n684), .ZN(G288) );
  AND2_X1 U776 ( .A1(n691), .A2(n686), .ZN(n687) );
  XNOR2_X1 U777 ( .A(KEYINPUT83), .B(n687), .ZN(n698) );
  XOR2_X1 U778 ( .A(G303), .B(KEYINPUT19), .Z(n689) );
  XOR2_X1 U779 ( .A(G290), .B(G299), .Z(n688) );
  XNOR2_X1 U780 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U781 ( .A(n690), .B(G305), .ZN(n692) );
  XNOR2_X1 U782 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n693), .B(G288), .ZN(n916) );
  XOR2_X1 U784 ( .A(n916), .B(n694), .Z(n695) );
  NAND2_X1 U785 ( .A1(n695), .A2(G868), .ZN(n696) );
  XNOR2_X1 U786 ( .A(KEYINPUT82), .B(n696), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(G295) );
  NAND2_X1 U788 ( .A1(G2084), .A2(G2078), .ZN(n699) );
  XOR2_X1 U789 ( .A(KEYINPUT20), .B(n699), .Z(n700) );
  NAND2_X1 U790 ( .A1(G2090), .A2(n700), .ZN(n701) );
  XNOR2_X1 U791 ( .A(KEYINPUT21), .B(n701), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n702), .A2(G2072), .ZN(G158) );
  NAND2_X1 U793 ( .A1(G69), .A2(G120), .ZN(n703) );
  NOR2_X1 U794 ( .A1(G237), .A2(n703), .ZN(n704) );
  NAND2_X1 U795 ( .A1(G108), .A2(n704), .ZN(n853) );
  NAND2_X1 U796 ( .A1(G567), .A2(n853), .ZN(n705) );
  XNOR2_X1 U797 ( .A(n705), .B(KEYINPUT85), .ZN(n711) );
  XOR2_X1 U798 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n707) );
  NAND2_X1 U799 ( .A1(G132), .A2(G82), .ZN(n706) );
  XNOR2_X1 U800 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n708), .A2(G96), .ZN(n709) );
  OR2_X1 U802 ( .A1(G218), .A2(n709), .ZN(n854) );
  AND2_X1 U803 ( .A1(G2106), .A2(n854), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n710), .ZN(G319) );
  INV_X1 U805 ( .A(G319), .ZN(n713) );
  NAND2_X1 U806 ( .A1(G661), .A2(G483), .ZN(n712) );
  NOR2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U808 ( .A(KEYINPUT86), .B(n714), .ZN(n848) );
  NAND2_X1 U809 ( .A1(G36), .A2(n848), .ZN(G176) );
  XNOR2_X1 U810 ( .A(KEYINPUT91), .B(n802), .ZN(n715) );
  INV_X1 U811 ( .A(n731), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n716), .A2(G1996), .ZN(n718) );
  INV_X1 U813 ( .A(KEYINPUT26), .ZN(n717) );
  XNOR2_X1 U814 ( .A(n718), .B(n717), .ZN(n721) );
  AND2_X1 U815 ( .A1(n731), .A2(G1341), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n727), .A2(n991), .ZN(n726) );
  INV_X1 U817 ( .A(G2067), .ZN(n868) );
  XNOR2_X1 U818 ( .A(n722), .B(KEYINPUT99), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n763), .A2(G1348), .ZN(n723) );
  NAND2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U823 ( .A(n730), .B(KEYINPUT100), .ZN(n740) );
  INV_X1 U824 ( .A(G2072), .ZN(n939) );
  NOR2_X1 U825 ( .A1(n731), .A2(n939), .ZN(n734) );
  XOR2_X1 U826 ( .A(KEYINPUT96), .B(KEYINPUT27), .Z(n732) );
  XNOR2_X1 U827 ( .A(KEYINPUT95), .B(n732), .ZN(n733) );
  XNOR2_X1 U828 ( .A(n734), .B(n733), .ZN(n736) );
  XOR2_X1 U829 ( .A(G1956), .B(KEYINPUT97), .Z(n1025) );
  NAND2_X1 U830 ( .A1(n763), .A2(n1025), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n994), .A2(n741), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n745) );
  NOR2_X1 U834 ( .A1(n741), .A2(n994), .ZN(n743) );
  INV_X1 U835 ( .A(KEYINPUT28), .ZN(n742) );
  XNOR2_X1 U836 ( .A(n743), .B(n742), .ZN(n744) );
  NAND2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U838 ( .A(KEYINPUT29), .B(n746), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n763), .A2(G1961), .ZN(n749) );
  XOR2_X1 U840 ( .A(G2078), .B(KEYINPUT25), .Z(n747) );
  XNOR2_X1 U841 ( .A(KEYINPUT92), .B(n747), .ZN(n973) );
  NAND2_X1 U842 ( .A1(n716), .A2(n973), .ZN(n748) );
  NAND2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U844 ( .A(n750), .B(KEYINPUT93), .ZN(n755) );
  NAND2_X1 U845 ( .A1(G171), .A2(n755), .ZN(n751) );
  XOR2_X1 U846 ( .A(KEYINPUT94), .B(n751), .Z(n752) );
  NOR2_X1 U847 ( .A1(n753), .A2(n752), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G8), .A2(n763), .ZN(n798) );
  NOR2_X1 U849 ( .A1(G2084), .A2(n763), .ZN(n772) );
  NOR2_X1 U850 ( .A1(G168), .A2(n754), .ZN(n757) );
  NOR2_X1 U851 ( .A1(G171), .A2(n755), .ZN(n756) );
  NOR2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U853 ( .A(n758), .B(KEYINPUT31), .ZN(n759) );
  NOR2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U855 ( .A(n761), .B(KEYINPUT101), .ZN(n774) );
  AND2_X1 U856 ( .A1(G286), .A2(G8), .ZN(n762) );
  NAND2_X1 U857 ( .A1(n774), .A2(n762), .ZN(n770) );
  NOR2_X1 U858 ( .A1(G1971), .A2(n798), .ZN(n765) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n763), .ZN(n764) );
  NOR2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U861 ( .A(KEYINPUT103), .B(n766), .Z(n767) );
  NAND2_X1 U862 ( .A1(n767), .A2(G303), .ZN(n768) );
  OR2_X1 U863 ( .A1(n541), .A2(n768), .ZN(n769) );
  NAND2_X1 U864 ( .A1(G8), .A2(n772), .ZN(n778) );
  INV_X1 U865 ( .A(KEYINPUT102), .ZN(n773) );
  XNOR2_X1 U866 ( .A(n774), .B(n773), .ZN(n775) );
  NOR2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U869 ( .A1(G1971), .A2(G303), .ZN(n781) );
  XOR2_X1 U870 ( .A(n781), .B(KEYINPUT104), .Z(n783) );
  NOR2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n999) );
  INV_X1 U872 ( .A(n999), .ZN(n782) );
  AND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n792), .A2(n784), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n997) );
  AND2_X1 U876 ( .A1(n997), .A2(n536), .ZN(n785) );
  XOR2_X1 U877 ( .A(G1981), .B(G305), .Z(n1007) );
  NAND2_X1 U878 ( .A1(n999), .A2(KEYINPUT33), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n798), .A2(n787), .ZN(n788) );
  NOR2_X1 U880 ( .A1(G2090), .A2(G303), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G8), .A2(n793), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n792), .A2(n794), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n798), .A2(n795), .ZN(n800) );
  NOR2_X1 U884 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U885 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  OR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n844) );
  XNOR2_X1 U888 ( .A(G1986), .B(G290), .ZN(n1003) );
  AND2_X1 U889 ( .A1(n844), .A2(n1003), .ZN(n831) );
  NAND2_X1 U890 ( .A1(G129), .A2(n899), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G141), .A2(n638), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n808) );
  NAND2_X1 U893 ( .A1(n902), .A2(G105), .ZN(n806) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n806), .Z(n807) );
  NOR2_X1 U895 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n898), .A2(G117), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n908) );
  NAND2_X1 U898 ( .A1(G1996), .A2(n908), .ZN(n818) );
  NAND2_X1 U899 ( .A1(G119), .A2(n899), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G95), .A2(n902), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n816) );
  NAND2_X1 U902 ( .A1(G107), .A2(n898), .ZN(n814) );
  NAND2_X1 U903 ( .A1(G131), .A2(n638), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n883) );
  NAND2_X1 U906 ( .A1(G1991), .A2(n883), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n947) );
  AND2_X1 U908 ( .A1(n844), .A2(n947), .ZN(n836) );
  XNOR2_X1 U909 ( .A(KEYINPUT89), .B(n836), .ZN(n828) );
  XOR2_X1 U910 ( .A(n868), .B(KEYINPUT37), .Z(n841) );
  NAND2_X1 U911 ( .A1(G104), .A2(n902), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G140), .A2(n638), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U914 ( .A(KEYINPUT34), .B(n821), .ZN(n826) );
  NAND2_X1 U915 ( .A1(G116), .A2(n898), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G128), .A2(n899), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT35), .B(n824), .Z(n825) );
  NOR2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U920 ( .A(KEYINPUT36), .B(n827), .ZN(n895) );
  NOR2_X1 U921 ( .A1(n841), .A2(n895), .ZN(n954) );
  NAND2_X1 U922 ( .A1(n844), .A2(n954), .ZN(n839) );
  NAND2_X1 U923 ( .A1(n828), .A2(n839), .ZN(n829) );
  XNOR2_X1 U924 ( .A(KEYINPUT90), .B(n829), .ZN(n830) );
  NOR2_X1 U925 ( .A1(G1996), .A2(n908), .ZN(n945) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n833) );
  NOR2_X1 U927 ( .A1(G1991), .A2(n883), .ZN(n832) );
  XOR2_X1 U928 ( .A(KEYINPUT107), .B(n832), .Z(n950) );
  NOR2_X1 U929 ( .A1(n833), .A2(n950), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n834), .B(KEYINPUT108), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U932 ( .A1(n945), .A2(n837), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n838), .B(KEYINPUT39), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n842) );
  NAND2_X1 U935 ( .A1(n841), .A2(n895), .ZN(n961) );
  NAND2_X1 U936 ( .A1(n842), .A2(n961), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n846), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n937), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U941 ( .A1(G661), .A2(n847), .ZN(G259) );
  INV_X1 U942 ( .A(n848), .ZN(n851) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n849) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(n849), .Z(n850) );
  NOR2_X1 U945 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U946 ( .A(KEYINPUT111), .B(n852), .ZN(G188) );
  INV_X1 U948 ( .A(G132), .ZN(G219) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G82), .ZN(G220) );
  INV_X1 U952 ( .A(G69), .ZN(G235) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U955 ( .A(G1996), .B(KEYINPUT41), .ZN(n864) );
  XOR2_X1 U956 ( .A(G1981), .B(G1956), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1991), .B(G1966), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1961), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U962 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U963 ( .A(KEYINPUT112), .B(G2474), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(G229) );
  XNOR2_X1 U966 ( .A(n865), .B(G2096), .ZN(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n872) );
  XOR2_X1 U969 ( .A(G2678), .B(G2090), .Z(n870) );
  XOR2_X1 U970 ( .A(n868), .B(G2072), .Z(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U972 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U973 ( .A(G2084), .B(G2078), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(G227) );
  NAND2_X1 U975 ( .A1(G136), .A2(n638), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G112), .A2(n898), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G100), .A2(n902), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n899), .A2(G124), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT44), .B(n877), .Z(n878) );
  NOR2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n882), .B(KEYINPUT113), .ZN(G162) );
  XNOR2_X1 U984 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n883), .B(G162), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n948), .B(n886), .ZN(n897) );
  NAND2_X1 U988 ( .A1(G115), .A2(n898), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G127), .A2(n899), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G103), .A2(n902), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n638), .A2(G139), .ZN(n892) );
  XOR2_X1 U995 ( .A(KEYINPUT114), .B(n892), .Z(n893) );
  NOR2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n938) );
  XNOR2_X1 U997 ( .A(n895), .B(n938), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n913) );
  NAND2_X1 U999 ( .A1(G118), .A2(n898), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G130), .A2(n899), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n902), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n638), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n905), .B(KEYINPUT45), .Z(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(G164), .B(n911), .Z(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G395) );
  INV_X1 U1011 ( .A(G171), .ZN(G301) );
  XOR2_X1 U1012 ( .A(G301), .B(G286), .Z(n919) );
  XOR2_X1 U1013 ( .A(n916), .B(n915), .Z(n917) );
  XNOR2_X1 U1014 ( .A(n917), .B(n1012), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n920), .ZN(G397) );
  XOR2_X1 U1017 ( .A(G2454), .B(G2430), .Z(n922) );
  XNOR2_X1 U1018 ( .A(G2451), .B(G2446), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n922), .B(n921), .ZN(n929) );
  XOR2_X1 U1020 ( .A(G2443), .B(G2427), .Z(n924) );
  XNOR2_X1 U1021 ( .A(G2438), .B(KEYINPUT109), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1023 ( .A(n925), .B(G2435), .Z(n927) );
  XNOR2_X1 U1024 ( .A(G1341), .B(G1348), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n927), .B(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n929), .B(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n930), .A2(G14), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(G319), .A2(n936), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(G229), .A2(G227), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(KEYINPUT49), .B(n931), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1034 ( .A(G225), .ZN(G308) );
  INV_X1 U1035 ( .A(G108), .ZN(G238) );
  INV_X1 U1036 ( .A(n936), .ZN(G401) );
  INV_X1 U1037 ( .A(n937), .ZN(G223) );
  XOR2_X1 U1038 ( .A(n939), .B(n938), .Z(n942) );
  XNOR2_X1 U1039 ( .A(G164), .B(G2078), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(KEYINPUT116), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(n943), .B(KEYINPUT50), .ZN(n959) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1045 ( .A(KEYINPUT51), .B(n946), .Z(n956) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1051 ( .A(KEYINPUT115), .B(n957), .Z(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n962), .B(KEYINPUT52), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT117), .B(n963), .ZN(n965) );
  INV_X1 U1056 ( .A(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n966), .A2(G29), .ZN(n1049) );
  XOR2_X1 U1059 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n980) );
  XOR2_X1 U1060 ( .A(G2072), .B(G33), .Z(n968) );
  XOR2_X1 U1061 ( .A(G2067), .B(G26), .Z(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1063 ( .A(G1991), .B(G25), .Z(n969) );
  NAND2_X1 U1064 ( .A1(n969), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT118), .B(n970), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(n973), .B(G27), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G32), .B(G1996), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1070 ( .A(KEYINPUT119), .B(n976), .Z(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n980), .B(n979), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G35), .B(G2090), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1075 ( .A(G2084), .B(G34), .Z(n983) );
  XNOR2_X1 U1076 ( .A(KEYINPUT54), .B(n983), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT55), .B(n986), .Z(n988) );
  INV_X1 U1079 ( .A(G29), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n989), .ZN(n1047) );
  XNOR2_X1 U1082 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n990) );
  XOR2_X1 U1083 ( .A(G16), .B(n990), .Z(n1018) );
  XOR2_X1 U1084 ( .A(G171), .B(G1961), .Z(n993) );
  XOR2_X1 U1085 ( .A(n991), .B(G1348), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1005) );
  XOR2_X1 U1087 ( .A(n994), .B(G1956), .Z(n996) );
  XOR2_X1 U1088 ( .A(G166), .B(G1971), .Z(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(KEYINPUT122), .B(n1001), .Z(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT123), .B(n1006), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT57), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(G1341), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT124), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1045) );
  INV_X1 U1105 ( .A(G16), .ZN(n1043) );
  XOR2_X1 U1106 ( .A(G1976), .B(G23), .Z(n1020) );
  XOR2_X1 U1107 ( .A(G1971), .B(G22), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(G24), .B(G1986), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1023), .Z(n1040) );
  XOR2_X1 U1112 ( .A(G1961), .B(G5), .Z(n1035) );
  XNOR2_X1 U1113 ( .A(G1348), .B(KEYINPUT59), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(n1024), .B(G4), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(n1025), .B(G20), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(G6), .B(G1981), .ZN(n1026) );
  NOR2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT126), .B(G1341), .ZN(n1030) );
  XNOR2_X1 U1120 ( .A(G19), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1122 ( .A(KEYINPUT60), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1123 ( .A1(n1035), .A2(n1034), .ZN(n1037) );
  XNOR2_X1 U1124 ( .A(G21), .B(G1966), .ZN(n1036) );
  NOR2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1126 ( .A(KEYINPUT127), .B(n1038), .ZN(n1039) );
  NOR2_X1 U1127 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1128 ( .A(KEYINPUT61), .B(n1041), .ZN(n1042) );
  NAND2_X1 U1129 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1130 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NOR2_X1 U1131 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NAND2_X1 U1132 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1133 ( .A(KEYINPUT62), .B(n1050), .ZN(G150) );
  INV_X1 U1134 ( .A(G150), .ZN(G311) );
endmodule

