//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(G567), .A2(new_n455), .B1(new_n452), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n459), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  INV_X1    g044(.A(new_n461), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n459), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n459), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n459), .ZN(new_n478));
  OAI221_X1 g053(.A(new_n473), .B1(new_n474), .B2(new_n475), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n482));
  OR2_X1    g057(.A1(G102), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n460), .B2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n461), .C2(new_n460), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  OR2_X1    g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT5), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(G166));
  XOR2_X1   g082(.A(KEYINPUT71), .B(G89), .Z(new_n508));
  INV_X1    g083(.A(G51), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n502), .A2(new_n508), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n510), .A2(new_n514), .ZN(G286));
  INV_X1    g090(.A(G286), .ZN(G168));
  NAND3_X1  g091(.A1(new_n501), .A2(G52), .A3(G543), .ZN(new_n517));
  INV_X1    g092(.A(G90), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n502), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n517), .B(KEYINPUT73), .C1(new_n502), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G77), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G64), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT72), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n532), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n523), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n535), .B1(new_n523), .B2(new_n534), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n499), .ZN(new_n540));
  OR2_X1    g115(.A1(KEYINPUT6), .A2(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(KEYINPUT6), .A2(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n495), .A2(new_n496), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n543), .A2(G81), .B1(new_n545), .B2(G43), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n495), .B2(new_n496), .ZN(new_n554));
  AND2_X1   g129(.A1(G78), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n543), .A2(G91), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n545), .B2(G53), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT6), .A2(G651), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT6), .A2(G651), .ZN(new_n561));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n556), .B(new_n557), .C1(new_n559), .C2(new_n563), .ZN(G299));
  NOR2_X1   g139(.A1(new_n536), .A2(new_n537), .ZN(G301));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n543), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n545), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n567), .A2(new_n572), .A3(new_n568), .A4(new_n569), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n497), .A2(new_n501), .A3(G86), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT77), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT76), .B1(new_n527), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n497), .A2(new_n580), .A3(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  AND2_X1   g160(.A1(G48), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(new_n501), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n560), .C2(new_n561), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n577), .A2(new_n584), .A3(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n499), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n502), .A2(new_n594), .B1(new_n504), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n543), .A2(G92), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT10), .Z(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n527), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n545), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  MUX2_X1   g184(.A(new_n599), .B(new_n608), .S(new_n609), .Z(G284));
  MUX2_X1   g185(.A(new_n599), .B(new_n608), .S(new_n609), .Z(G321));
  XOR2_X1   g186(.A(G299), .B(KEYINPUT80), .Z(new_n612));
  MUX2_X1   g187(.A(new_n612), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g188(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n607), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n477), .A2(new_n466), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n472), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n459), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n478), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n638), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT84), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n656), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n657), .B(new_n659), .C1(new_n652), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n652), .A3(new_n655), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n659), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n664), .B1(new_n665), .B2(new_n654), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G1986), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n673), .A2(new_n674), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(new_n675), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n678), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n682), .B1(new_n681), .B2(new_n685), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n672), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(G1986), .A3(new_n686), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n671), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT89), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n689), .A2(new_n691), .A3(new_n671), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n696), .ZN(new_n699));
  INV_X1    g274(.A(new_n697), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G2090), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT100), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(G33), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT93), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(new_n459), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n715), .ZN(new_n719));
  INV_X1    g294(.A(G139), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n478), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n711), .B1(new_n722), .B2(new_n704), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2072), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n704), .A2(G32), .ZN(new_n725));
  INV_X1    g300(.A(new_n478), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n726), .A2(G141), .B1(G129), .B2(new_n472), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n728));
  AND3_X1   g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n730), .A2(new_n731), .B1(G105), .B2(new_n466), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n725), .B1(new_n734), .B2(new_n704), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT96), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n704), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G2084), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n724), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT97), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n710), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G171), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT98), .B(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n736), .A2(new_n737), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n607), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT90), .B(G1348), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n704), .A2(G26), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT28), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n472), .A2(G128), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT92), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n726), .A2(G140), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n459), .A2(G116), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  INV_X1    g341(.A(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G20), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  INV_X1    g344(.A(G299), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n767), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n752), .A2(new_n756), .A3(new_n766), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n767), .A2(G19), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n547), .B2(new_n767), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT91), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G28), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n704), .B1(new_n780), .B2(G28), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .C1(new_n631), .C2(new_n704), .ZN(new_n783));
  NOR2_X1   g358(.A1(G27), .A2(G29), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G164), .B2(G29), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n783), .B1(G2078), .B2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  INV_X1    g363(.A(new_n743), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n767), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n767), .ZN(new_n793));
  INV_X1    g368(.A(G1966), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n778), .A2(new_n786), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n774), .B(new_n796), .C1(G2090), .C2(new_n708), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n747), .A2(new_n751), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n767), .A2(G23), .ZN(new_n799));
  INV_X1    g374(.A(new_n570), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n767), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n767), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n767), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1971), .ZN(new_n806));
  INV_X1    g381(.A(G305), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G6), .B2(G16), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT32), .B(G1981), .Z(new_n810));
  AOI211_X1 g385(.A(new_n803), .B(new_n806), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n704), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n726), .A2(G131), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n472), .A2(G119), .ZN(new_n817));
  OR2_X1    g392(.A1(G95), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n704), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(G16), .A2(G24), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n597), .B2(G16), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1986), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n813), .A2(new_n814), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n798), .B1(new_n831), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n831), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n834), .A2(new_n751), .A3(new_n797), .A4(new_n747), .ZN(G150));
  AOI22_X1  g410(.A1(new_n497), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n499), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n502), .A2(new_n838), .B1(new_n504), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n606), .A2(new_n615), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n547), .B(new_n841), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n850), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(G145));
  XOR2_X1   g428(.A(new_n631), .B(G160), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n764), .B(G164), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n722), .A2(new_n734), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n733), .B1(new_n718), .B2(new_n721), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n821), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n821), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n857), .A3(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n472), .A2(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n459), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(G142), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n868), .B1(new_n869), .B2(new_n870), .C1(new_n871), .C2(new_n478), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n622), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n867), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n873), .B1(new_n865), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n856), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n879), .A2(new_n875), .A3(new_n855), .A4(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g458(.A(new_n597), .B(new_n800), .ZN(new_n884));
  OR2_X1    g459(.A1(G166), .A2(KEYINPUT103), .ZN(new_n885));
  NAND2_X1  g460(.A1(G166), .A2(KEYINPUT103), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n807), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(G305), .A3(new_n886), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n884), .A3(new_n889), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT42), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  INV_X1    g469(.A(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n893), .B1(new_n898), .B2(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n606), .B(new_n770), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n848), .B(new_n617), .ZN(new_n903));
  MUX2_X1   g478(.A(new_n900), .B(new_n902), .S(new_n903), .Z(new_n904));
  XOR2_X1   g479(.A(new_n899), .B(new_n904), .Z(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G868), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g482(.A(new_n906), .B1(G868), .B2(new_n841), .ZN(G331));
  XOR2_X1   g483(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n909));
  INV_X1    g484(.A(new_n848), .ZN(new_n910));
  NAND2_X1  g485(.A1(G301), .A2(G286), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(G301), .A2(G286), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(G171), .A2(G168), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n848), .A3(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n902), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n900), .A3(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n920), .B2(new_n898), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n918), .A2(new_n897), .A3(new_n896), .A4(new_n919), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n909), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n920), .A2(new_n898), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n923), .A3(new_n881), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT44), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(G397));
  NAND2_X1  g508(.A1(new_n491), .A2(new_n493), .ZN(new_n934));
  INV_X1    g509(.A(new_n487), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G40), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n464), .A2(new_n468), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(KEYINPUT111), .B(G8), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT49), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n576), .B1(new_n587), .B2(new_n589), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n949), .B1(new_n583), .B2(G651), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT113), .B(new_n576), .C1(new_n587), .C2(new_n589), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n682), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n577), .A2(new_n584), .A3(new_n682), .A4(new_n590), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n949), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n956), .A2(new_n584), .A3(new_n951), .ZN(new_n957));
  OAI211_X1 g532(.A(KEYINPUT49), .B(new_n953), .C1(new_n957), .C2(new_n682), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n946), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n800), .A2(G1976), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n944), .B1(new_n939), .B2(new_n941), .ZN(new_n961));
  AOI211_X1 g536(.A(KEYINPUT112), .B(new_n940), .C1(new_n936), .C2(new_n938), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT52), .ZN(new_n964));
  INV_X1    g539(.A(G1976), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n571), .A2(new_n965), .A3(new_n573), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(new_n960), .C1(new_n962), .C2(new_n961), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n959), .A2(new_n964), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT109), .B(G1971), .Z(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1384), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n938), .B1(G164), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n493), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n492), .B1(new_n477), .B2(new_n489), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n482), .B(new_n486), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n972), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n983));
  INV_X1    g558(.A(G2090), .ZN(new_n984));
  NOR2_X1   g559(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n983), .A2(new_n984), .A3(new_n938), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n971), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n500), .B2(new_n506), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n989), .B(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT110), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n982), .A2(new_n987), .ZN(new_n993));
  AND4_X1   g568(.A1(KEYINPUT110), .A2(new_n993), .A3(G8), .A4(new_n991), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n970), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n955), .A2(new_n958), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n574), .A2(new_n965), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n953), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n946), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(G286), .A2(new_n941), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n794), .B1(new_n976), .B2(new_n981), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n983), .A2(new_n790), .A3(new_n938), .A4(new_n986), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n971), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1000), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT51), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n940), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n1009), .B2(new_n1000), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT120), .A3(new_n1007), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n994), .A2(new_n992), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n991), .B1(new_n993), .B2(new_n941), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n970), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n973), .B1(G164), .B2(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n979), .A2(new_n974), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n788), .A3(new_n938), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1961), .ZN(new_n1030));
  INV_X1    g605(.A(new_n985), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n938), .B1(G164), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n979), .B2(new_n980), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1028), .A2(G2078), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1025), .A2(new_n938), .A3(new_n1026), .A4(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1029), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G171), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1024), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n999), .B1(new_n1021), .B2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1009), .A2(G286), .A3(new_n940), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1024), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT63), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1022), .A2(new_n970), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n988), .A2(new_n991), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1043), .A2(new_n1047), .A3(KEYINPUT63), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1044), .A2(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT107), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n936), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT107), .B1(G164), .B2(G1384), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n973), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n462), .A2(new_n463), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n459), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  NOR4_X1   g633(.A1(new_n468), .A2(new_n1028), .A3(new_n937), .A4(G2078), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1054), .A2(new_n1026), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(G301), .A3(new_n1029), .A4(new_n1035), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1039), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1011), .A2(new_n1016), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G171), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1038), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1063), .B1(new_n1069), .B2(G301), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1024), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1024), .A2(new_n1064), .A3(KEYINPUT124), .A4(new_n1072), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n1077));
  AND3_X1   g652(.A1(G299), .A2(new_n1077), .A3(KEYINPUT57), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(G299), .B2(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n772), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1025), .A2(new_n938), .A3(new_n1026), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1081), .A2(KEYINPUT115), .A3(new_n1083), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1080), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n939), .ZN(new_n1090));
  INV_X1    g665(.A(G2067), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(G1348), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n607), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1085), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1025), .A2(new_n938), .A3(new_n1026), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT58), .B(G1341), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1097), .A2(G1996), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n547), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1084), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1080), .A2(new_n1081), .A3(KEYINPUT117), .A4(new_n1083), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT61), .B1(new_n1088), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1080), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT116), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1084), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1102), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1092), .B(KEYINPUT60), .C1(new_n1093), .C2(G1348), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1117), .A2(KEYINPUT118), .A3(new_n606), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n606), .B1(new_n1117), .B2(KEYINPUT118), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(KEYINPUT118), .B2(new_n1117), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1094), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(KEYINPUT60), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1096), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1075), .B(new_n1076), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1050), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(G160), .A2(G40), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1054), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n764), .B(new_n1091), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n733), .A2(G1996), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n733), .A2(G1996), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1130), .A2(KEYINPUT108), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT108), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n821), .A2(new_n823), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n820), .A2(new_n824), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1129), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n597), .B(new_n672), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1129), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1127), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1130), .A2(G1996), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT46), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1130), .B1(new_n1131), .B2(new_n734), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT47), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(G2067), .B2(new_n764), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1129), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT125), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1129), .A2(new_n672), .A3(new_n597), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT48), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1137), .A2(new_n1158), .A3(new_n1140), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1155), .A2(KEYINPUT125), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1144), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1165));
  OAI21_X1  g739(.A(G319), .B1(new_n649), .B2(new_n650), .ZN(new_n1166));
  NOR2_X1   g740(.A1(G227), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g741(.A1(new_n702), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n702), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g743(.A(new_n882), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n924), .A2(new_n925), .ZN(new_n1171));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n1171), .ZN(G308));
  OAI221_X1 g746(.A(new_n882), .B1(new_n924), .B2(new_n925), .C1(new_n1169), .C2(new_n1168), .ZN(G225));
endmodule


