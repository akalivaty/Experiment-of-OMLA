//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  INV_X1    g026(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n452), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g052(.A(KEYINPUT69), .B(G2105), .C1(new_n469), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(G137), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G101), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(new_n481), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n495), .B2(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n494), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n492), .B2(new_n493), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n502), .B(new_n505), .C1(new_n493), .C2(new_n492), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(G126), .B(G2105), .C1(new_n492), .C2(new_n493), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n481), .A2(G114), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n508), .B(KEYINPUT70), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n467), .B2(new_n468), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n507), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  OR2_X1    g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n528), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n524), .A2(new_n534), .ZN(G166));
  INV_X1    g110(.A(new_n521), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n531), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n529), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(new_n529), .A2(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n532), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n521), .A2(G64), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n523), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n521), .A2(G56), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n523), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(KEYINPUT71), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n556));
  AOI211_X1 g131(.A(new_n556), .B(new_n523), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n529), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n532), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g135(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT72), .Z(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT73), .Z(G188));
  NAND2_X1  g143(.A1(new_n529), .A2(G53), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n536), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n519), .A2(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n573), .A2(G651), .B1(G91), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(new_n547), .B2(new_n550), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n574), .A2(G90), .B1(new_n529), .B2(G52), .ZN(new_n579));
  INV_X1    g154(.A(G64), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n519), .B2(new_n520), .ZN(new_n581));
  INV_X1    g156(.A(new_n549), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n579), .A2(KEYINPUT74), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G301));
  INV_X1    g161(.A(G168), .ZN(G286));
  OR2_X1    g162(.A1(new_n524), .A2(new_n534), .ZN(G303));
  OAI21_X1  g163(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n529), .A2(G49), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n532), .ZN(G288));
  NAND2_X1  g167(.A1(new_n574), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n529), .A2(G48), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n523), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n595), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n523), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n529), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n532), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n600), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n536), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n532), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n574), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT75), .B1(new_n615), .B2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n585), .A2(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n616), .B(KEYINPUT75), .S(new_n618), .Z(G284));
  XNOR2_X1  g194(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n615), .B1(new_n625), .B2(G860), .ZN(G148));
  OR3_X1    g201(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n617), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n614), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n617), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n480), .A2(new_n484), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XOR2_X1   g208(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n495), .A2(G123), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT78), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(G111), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G2105), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n497), .B2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n636), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(G2096), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n637), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT80), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G1341), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G1348), .ZN(new_n664));
  INV_X1    g239(.A(G1341), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G1348), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n654), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G14), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n668), .A3(new_n654), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  INV_X1    g253(.A(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n674), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n676), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n683), .B2(new_n679), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n679), .A3(new_n674), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n690), .A2(new_n695), .A3(new_n693), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n698));
  AOI211_X1 g273(.A(new_n694), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1981), .B(G1986), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n700), .B(new_n701), .ZN(new_n709));
  INV_X1    g284(.A(new_n707), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(G229));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT86), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n497), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n495), .A2(G119), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n481), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G24), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n600), .A2(new_n603), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1986), .Z(new_n728));
  OR2_X1    g303(.A1(G16), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n730));
  OR2_X1    g305(.A1(G288), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G288), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n729), .B1(new_n733), .B2(new_n724), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT33), .B(G1976), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n724), .A2(G22), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G166), .B2(new_n724), .ZN(new_n739));
  INV_X1    g314(.A(G1971), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G6), .A2(G16), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n595), .A2(new_n597), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G16), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT32), .B(G1981), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n736), .A2(new_n737), .A3(new_n741), .A4(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n723), .B(new_n728), .C1(new_n747), .C2(KEYINPUT34), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(KEYINPUT34), .B2(new_n747), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  NOR2_X1   g328(.A1(G168), .A2(new_n724), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n724), .B2(G21), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n480), .A2(new_n481), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(new_n481), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n713), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n713), .B2(G33), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n757), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n758), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n724), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n724), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1961), .ZN(new_n774));
  INV_X1    g349(.A(G11), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT31), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT31), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n713), .B1(new_n778), .B2(G28), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n777), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n644), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G29), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n495), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n484), .A2(G105), .ZN(new_n788));
  INV_X1    g363(.A(G141), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n763), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n713), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n713), .B2(G32), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n783), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n771), .A2(new_n774), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT93), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n713), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n713), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2078), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n713), .A2(G26), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT28), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n480), .A2(G140), .A3(new_n481), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n480), .A2(G128), .A3(G2105), .ZN(new_n806));
  OR2_X1    g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G116), .C2(new_n481), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT89), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(KEYINPUT89), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n724), .A2(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n561), .B2(new_n724), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n665), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n796), .A2(new_n802), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n724), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT23), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n622), .B2(new_n724), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1956), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n713), .A2(G35), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G162), .B2(new_n713), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT29), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n823), .B1(new_n827), .B2(G2090), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n724), .A2(G4), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n615), .B2(new_n724), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1348), .ZN(new_n833));
  INV_X1    g408(.A(G2084), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n835));
  AOI21_X1  g410(.A(G29), .B1(new_n835), .B2(G34), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G34), .B2(new_n835), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT91), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n487), .B2(new_n713), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n833), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n755), .A2(new_n756), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT94), .ZN(new_n842));
  INV_X1    g417(.A(G2090), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n826), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n830), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n839), .A2(new_n834), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT92), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n828), .B2(new_n829), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n819), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n752), .A2(new_n753), .A3(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI211_X1 g428(.A(KEYINPUT96), .B(new_n852), .C1(new_n536), .C2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n853), .B1(new_n519), .B2(new_n520), .ZN(new_n856));
  INV_X1    g431(.A(new_n852), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(G651), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n574), .A2(G93), .B1(new_n529), .B2(G55), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(KEYINPUT97), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT97), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n627), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n561), .A2(new_n859), .A3(new_n860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT38), .Z(new_n867));
  NOR2_X1   g442(.A1(new_n614), .A2(new_n625), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g447(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  NAND2_X1  g450(.A1(new_n497), .A2(G142), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n495), .A2(G130), .ZN(new_n877));
  OR2_X1    g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G2104), .C1(G118), .C2(new_n481), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT103), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(new_n633), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n880), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n633), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n720), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n881), .A2(new_n633), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n885), .ZN(new_n889));
  INV_X1    g464(.A(new_n720), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n494), .A2(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n504), .B2(new_n506), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n809), .ZN(new_n895));
  INV_X1    g470(.A(new_n809), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n514), .A2(new_n515), .ZN(new_n897));
  INV_X1    g472(.A(new_n506), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n505), .B1(new_n480), .B2(new_n502), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n791), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n791), .A2(new_n895), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT100), .ZN(new_n907));
  INV_X1    g482(.A(new_n767), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n906), .B2(KEYINPUT100), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n911));
  INV_X1    g486(.A(new_n905), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n791), .B1(new_n895), .B2(new_n901), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT101), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n904), .A2(new_n915), .A3(new_n905), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n917), .B2(new_n908), .ZN(new_n918));
  AOI211_X1 g493(.A(KEYINPUT102), .B(new_n767), .C1(new_n914), .C2(new_n916), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n892), .B(new_n910), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n910), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(new_n892), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n644), .B(new_n499), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(G160), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(G160), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n933), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n937), .A2(new_n920), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n940), .B2(new_n925), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g518(.A1(new_n733), .A2(new_n743), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G166), .ZN(new_n945));
  NAND2_X1  g520(.A1(G303), .A2(new_n726), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G305), .B1(new_n731), .B2(new_n732), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n944), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  OR3_X1    g530(.A1(new_n951), .A2(new_n955), .A3(KEYINPUT42), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n951), .B2(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n866), .B(new_n629), .ZN(new_n960));
  NAND2_X1  g535(.A1(G299), .A2(new_n614), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n570), .A2(new_n575), .A3(new_n608), .A4(new_n613), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n961), .A2(KEYINPUT41), .A3(new_n962), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT41), .B1(new_n961), .B2(new_n962), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n969), .B2(new_n960), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n617), .B1(new_n959), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n954), .A2(new_n958), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT107), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n617), .B1(new_n862), .B2(new_n863), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n972), .B2(new_n974), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n976), .A2(new_n979), .ZN(G295));
  NOR2_X1   g555(.A1(new_n976), .A2(new_n979), .ZN(G331));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n951), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT109), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n859), .A2(new_n860), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT97), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n561), .B1(new_n988), .B2(new_n861), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n627), .A2(new_n986), .ZN(new_n990));
  NOR2_X1   g565(.A1(G171), .A2(G168), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n585), .B2(G168), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n547), .A2(new_n550), .A3(new_n577), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT74), .B1(new_n579), .B2(new_n583), .ZN(new_n995));
  OAI21_X1  g570(.A(G168), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G168), .B2(G171), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n864), .B2(new_n865), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n964), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n989), .B2(new_n990), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n864), .A3(new_n865), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n968), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT108), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(KEYINPUT108), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n985), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n968), .A2(new_n1001), .A3(new_n1000), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n963), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n951), .A3(new_n1004), .ZN(new_n1011));
  INV_X1    g586(.A(G37), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1006), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT43), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n999), .A2(new_n1002), .ZN(new_n1015));
  AOI21_X1  g590(.A(G37), .B1(new_n985), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1011), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(KEYINPUT44), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n1012), .A3(new_n1006), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1026), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n900), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n486), .A2(new_n1031), .A3(G40), .A4(new_n475), .ZN(new_n1032));
  INV_X1    g607(.A(new_n474), .ZN(new_n1033));
  OAI21_X1  g608(.A(G125), .B1(new_n492), .B2(new_n493), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n481), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n482), .A2(G40), .A3(new_n485), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT120), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1030), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G2078), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1039), .A2(KEYINPUT53), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n507), .B2(new_n897), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n517), .A2(new_n1029), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n477), .B2(new_n478), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n900), .A2(new_n1047), .A3(new_n1029), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT114), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1041), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1045), .A2(new_n1046), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1961), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1044), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT113), .A3(new_n1046), .A4(new_n1030), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1046), .A2(new_n1030), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT45), .B1(new_n517), .B2(new_n1029), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G2078), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(G301), .B(new_n1054), .C1(new_n1062), .C2(KEYINPUT53), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n517), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1055), .B1(new_n894), .B2(G1384), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1046), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1052), .A2(new_n1053), .B1(new_n1069), .B2(new_n1040), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1062), .B2(KEYINPUT53), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1064), .A2(new_n1065), .B1(new_n585), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1063), .A2(KEYINPUT121), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT54), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1057), .A2(new_n1061), .A3(new_n740), .ZN(new_n1075));
  AOI211_X1 g650(.A(G2090), .B(new_n1036), .C1(new_n477), .C2(new_n478), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1045), .A2(new_n1049), .A3(new_n1076), .A4(new_n1051), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT115), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n894), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1079), .A2(new_n1050), .B1(new_n1044), .B2(KEYINPUT50), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1049), .A4(new_n1076), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1075), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G303), .A2(G8), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT55), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(G8), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  INV_X1    g663(.A(G1981), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n743), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n743), .A2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT49), .A3(new_n1090), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1046), .A2(new_n1041), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(G8), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n731), .A2(G1976), .A3(new_n732), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(G8), .A3(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT52), .ZN(new_n1101));
  INV_X1    g676(.A(G1976), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(G288), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1097), .A2(new_n1099), .A3(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1098), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1087), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n1107), .B2(new_n1039), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1054), .ZN(new_n1109));
  OAI21_X1  g684(.A(G171), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1070), .B(G301), .C1(new_n1062), .C2(KEYINPUT53), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(KEYINPUT54), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT50), .B1(new_n894), .B2(G1384), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1046), .C1(new_n1044), .C2(KEYINPUT50), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1075), .B1(G2090), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G8), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1085), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1068), .A2(new_n756), .ZN(new_n1118));
  AOI211_X1 g693(.A(G2084), .B(new_n1036), .C1(new_n477), .C2(new_n478), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1045), .A2(new_n1049), .A3(new_n1119), .A4(new_n1051), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1120), .A3(G168), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G8), .ZN(new_n1122));
  AOI21_X1  g697(.A(G168), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT51), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1125), .A3(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1106), .A2(new_n1112), .A3(new_n1117), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1028), .B1(new_n1074), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1108), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(new_n1065), .A3(G301), .A4(new_n1054), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1071), .A2(new_n585), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1073), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1112), .A2(new_n1127), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1117), .A2(new_n1087), .A3(new_n1105), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT122), .A4(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(G299), .B(KEYINPUT57), .Z(new_n1139));
  INV_X1    g714(.A(G1956), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1114), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1056), .A2(new_n1046), .A3(new_n1030), .A4(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n614), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1096), .B(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n814), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1052), .A2(new_n667), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1139), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1144), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT58), .B(G1341), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1056), .A2(new_n1046), .A3(new_n1030), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1147), .A2(new_n1160), .B1(G1996), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(new_n561), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1139), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1157), .B1(new_n1144), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1162), .A2(new_n561), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(KEYINPUT119), .A3(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1159), .A2(new_n1164), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n615), .B1(new_n1150), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n614), .A4(new_n1149), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1172), .A2(new_n1173), .B1(new_n1171), .B2(new_n1150), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1156), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1129), .A2(new_n1138), .A3(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1127), .B(KEYINPUT62), .Z(new_n1177));
  NAND4_X1  g752(.A1(new_n1177), .A2(new_n585), .A3(new_n1137), .A4(new_n1071), .ZN(new_n1178));
  NAND2_X1  g753(.A1(G168), .A2(G8), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1117), .A2(new_n1087), .A3(new_n1105), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(KEYINPUT63), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1083), .A2(G8), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1184), .B2(new_n1085), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1181), .A2(new_n1182), .B1(new_n1185), .B2(new_n1106), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1105), .A2(G8), .A3(new_n1086), .A4(new_n1083), .ZN(new_n1187));
  NOR2_X1   g762(.A1(G288), .A2(G1976), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1098), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1097), .B1(new_n1189), .B2(new_n1091), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT116), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT116), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1191), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1106), .A2(new_n1185), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1193), .B(new_n1194), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1176), .A2(new_n1178), .A3(new_n1192), .A4(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1041), .A2(KEYINPUT45), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1046), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1200), .A2(G1996), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n791), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT111), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1200), .B(KEYINPUT112), .Z(new_n1204));
  NAND2_X1  g779(.A1(new_n896), .A2(new_n814), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n809), .A2(G2067), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(G1996), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1207), .B1(new_n1208), .B2(new_n791), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n720), .B(new_n722), .Z(new_n1212));
  NAND2_X1  g787(.A1(new_n1204), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1200), .ZN(new_n1215));
  XNOR2_X1  g790(.A(G290), .B(G1986), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1198), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1207), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1204), .B1(new_n903), .B2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1201), .B(KEYINPUT46), .Z(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(KEYINPUT123), .B(KEYINPUT47), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1214), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(KEYINPUT124), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1227));
  NOR3_X1   g802(.A1(new_n1200), .A2(G1986), .A3(G290), .ZN(new_n1228));
  XNOR2_X1  g803(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1229));
  XOR2_X1   g804(.A(new_n1228), .B(new_n1229), .Z(new_n1230));
  NOR3_X1   g805(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1211), .A2(new_n722), .A3(new_n890), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1205), .ZN(new_n1233));
  AOI211_X1 g808(.A(new_n1224), .B(new_n1231), .C1(new_n1204), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1218), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1237));
  NOR2_X1   g811(.A1(new_n464), .A2(G227), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n708), .A2(new_n711), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g813(.A(new_n1239), .B1(new_n671), .B2(new_n672), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n937), .B1(new_n926), .B2(new_n927), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n937), .A2(new_n920), .ZN(new_n1242));
  INV_X1    g816(.A(new_n925), .ZN(new_n1243));
  OAI21_X1  g817(.A(new_n1012), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g818(.A(new_n1240), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g819(.A1(new_n1016), .A2(new_n1024), .B1(new_n1013), .B2(KEYINPUT43), .ZN(new_n1246));
  OAI21_X1  g820(.A(new_n1237), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g821(.A1(new_n942), .A2(new_n1019), .A3(KEYINPUT126), .A4(new_n1240), .ZN(new_n1248));
  AND2_X1   g822(.A1(new_n1247), .A2(new_n1248), .ZN(G308));
  NAND2_X1  g823(.A1(new_n1247), .A2(new_n1248), .ZN(G225));
endmodule


