//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1251, new_n1252,
    new_n1253;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(G2104), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n458), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n471), .B(G2104), .C1(new_n461), .C2(new_n462), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n464), .A2(new_n465), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n460), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(new_n460), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G125), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT67), .A3(G125), .ZN(new_n486));
  NAND2_X1  g061(.A1(G113), .A2(G2104), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n476), .A2(new_n478), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n476), .A2(KEYINPUT72), .A3(new_n478), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(G160));
  NAND4_X1  g069(.A1(new_n464), .A2(G2105), .A3(new_n470), .A4(new_n472), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n497), .B(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G112), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n473), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G136), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(G162));
  INV_X1    g080(.A(G126), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n465), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n495), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n465), .A2(G138), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n485), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n464), .A2(new_n470), .A3(new_n472), .A4(new_n511), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT4), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G164));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n517), .A2(KEYINPUT6), .A3(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT6), .B1(new_n517), .B2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n522), .A2(G50), .B1(G651), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n518), .A2(new_n519), .ZN(new_n530));
  INV_X1    g105(.A(new_n526), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(KEYINPUT75), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n533), .B1(new_n520), .B2(new_n526), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G88), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n532), .A2(new_n534), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(G89), .ZN(G168));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT76), .B(G52), .Z(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n526), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n522), .A2(new_n549), .B1(new_n552), .B2(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND3_X1  g130(.A1(new_n532), .A2(G81), .A3(new_n534), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n526), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n522), .A2(G43), .B1(G651), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n556), .A2(new_n560), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n542), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n522), .B(G53), .C1(KEYINPUT79), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(G65), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(G65), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n531), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G78), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n521), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n532), .A2(G91), .A3(new_n534), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G299));
  INV_X1    g163(.A(G168), .ZN(G286));
  XNOR2_X1  g164(.A(new_n537), .B(KEYINPUT81), .ZN(G303));
  NAND2_X1  g165(.A1(new_n545), .A2(G87), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n531), .A2(G74), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n522), .B2(G49), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(new_n545), .A2(G86), .B1(G48), .B2(new_n522), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n526), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n595), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n545), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n526), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n522), .A2(G47), .B1(G651), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT83), .Z(new_n610));
  NAND3_X1  g185(.A1(new_n545), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n535), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT84), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n526), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(G651), .A2(new_n619), .B1(new_n522), .B2(G54), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n610), .B1(G868), .B2(new_n622), .ZN(G284));
  OAI21_X1  g198(.A(new_n610), .B1(G868), .B2(new_n622), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n587), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(G868), .B2(new_n587), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n634));
  NOR3_X1   g209(.A1(new_n467), .A2(new_n458), .A3(G2105), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n634), .B(new_n635), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2100), .Z(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n495), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G135), .B2(new_n503), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n638), .A2(new_n645), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT14), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n665), .B(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n674), .B2(new_n671), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n671), .A3(new_n668), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n670), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT92), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n692), .A2(new_n697), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n693), .A2(new_n697), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n685), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n698), .A3(new_n684), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n709), .B1(new_n705), .B2(new_n707), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n682), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n684), .B1(new_n706), .B2(new_n698), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n699), .A2(new_n704), .A3(new_n685), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n708), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n716), .A2(new_n681), .A3(new_n710), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G6), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n595), .A2(new_n601), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT95), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n719), .A2(G23), .ZN(new_n728));
  INV_X1    g303(.A(G288), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT33), .B(G1976), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n719), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n719), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1971), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n726), .A2(new_n727), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n726), .A2(new_n727), .A3(new_n739), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n740), .A3(KEYINPUT34), .ZN(new_n744));
  INV_X1    g319(.A(new_n495), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G119), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT93), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(G107), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n503), .B2(G131), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G25), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT35), .B(G1991), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT94), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n755), .A2(new_n757), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n719), .A2(G24), .ZN(new_n761));
  INV_X1    g336(.A(G290), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n719), .ZN(new_n763));
  INV_X1    g338(.A(G1986), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n759), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n743), .A2(new_n744), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(KEYINPUT36), .ZN(new_n769));
  INV_X1    g344(.A(new_n767), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n741), .B2(new_n742), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n771), .A2(new_n772), .A3(new_n744), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G160), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2084), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n719), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n719), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT102), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1966), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT103), .ZN(new_n783));
  INV_X1    g358(.A(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT30), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G29), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n719), .A2(G5), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G301), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1961), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n789), .B1(new_n790), .B2(new_n644), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G1966), .B2(new_n781), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n783), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(KEYINPUT104), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT104), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n783), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n778), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n719), .A2(G19), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n566), .B2(new_n719), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1341), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n719), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n622), .B2(new_n719), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n790), .A2(G32), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n503), .A2(G141), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT26), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n812), .A2(new_n813), .B1(G105), .B2(new_n459), .ZN(new_n814));
  INV_X1    g389(.A(G129), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n495), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n808), .B1(new_n817), .B2(new_n790), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT27), .B(G1996), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(new_n793), .B2(new_n792), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n803), .A2(new_n807), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n719), .A2(G20), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT23), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n587), .B2(new_n719), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1956), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n790), .A2(G26), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT28), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n472), .A2(new_n470), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT69), .B(KEYINPUT3), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n471), .B1(new_n830), .B2(G2104), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n832), .A2(KEYINPUT97), .A3(G128), .A4(G2105), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n834));
  INV_X1    g409(.A(G128), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n495), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G116), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G140), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n473), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n828), .B1(new_n845), .B2(G29), .ZN(new_n846));
  INV_X1    g421(.A(G2067), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(G27), .A2(G29), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G164), .B2(G29), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(G2078), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(G2078), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n819), .B2(new_n820), .ZN(new_n853));
  NOR4_X1   g428(.A1(new_n826), .A2(new_n848), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n822), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(G162), .A2(G29), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G29), .B2(G35), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT29), .ZN(new_n858));
  INV_X1    g433(.A(G2090), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n857), .A2(KEYINPUT29), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(KEYINPUT29), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(G2090), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(G29), .A2(G33), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT98), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT25), .Z(new_n868));
  INV_X1    g443(.A(G139), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n473), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(KEYINPUT99), .B(new_n868), .C1(new_n473), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(new_n465), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n866), .B1(new_n877), .B2(new_n790), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT100), .Z(new_n879));
  INV_X1    g454(.A(G2072), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n855), .A2(new_n864), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT101), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n800), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n800), .A2(new_n882), .A3(KEYINPUT105), .A4(new_n884), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n769), .A2(new_n773), .B1(new_n887), .B2(new_n888), .ZN(G311));
  NAND2_X1  g464(.A1(new_n769), .A2(new_n773), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(G150));
  NAND2_X1  g467(.A1(new_n562), .A2(new_n565), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n894));
  INV_X1    g469(.A(G651), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G55), .ZN(new_n897));
  INV_X1    g472(.A(G93), .ZN(new_n898));
  OAI221_X1 g473(.A(new_n896), .B1(new_n897), .B2(new_n542), .C1(new_n535), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n561), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n622), .A2(G559), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n907));
  AOI21_X1  g482(.A(G860), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(G860), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n910), .B(KEYINPUT37), .Z(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT106), .ZN(G145));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n914));
  INV_X1    g489(.A(new_n817), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n843), .B1(new_n836), .B2(new_n833), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n507), .A2(new_n508), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n745), .B2(G126), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n514), .A2(KEYINPUT4), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n512), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n509), .A2(new_n515), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT107), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n509), .B2(new_n515), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n845), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n924), .A2(new_n877), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n877), .B1(new_n924), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(G106), .A2(G2105), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n932));
  INV_X1    g507(.A(G130), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n495), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G142), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n473), .A2(new_n935), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT108), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT108), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n636), .ZN(new_n940));
  INV_X1    g515(.A(new_n636), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n753), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n942), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n937), .B2(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n752), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n877), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n921), .A2(new_n923), .A3(new_n916), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n845), .B1(new_n926), .B2(new_n925), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n924), .A2(new_n877), .A3(new_n927), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n817), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n930), .A2(new_n947), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G162), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n492), .A2(new_n493), .A3(new_n644), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n644), .B1(new_n492), .B2(new_n493), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G160), .A2(new_n643), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n492), .A2(new_n493), .A3(new_n644), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(G162), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n947), .B1(new_n930), .B2(new_n953), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n914), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n943), .A2(new_n946), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n928), .A2(new_n929), .A3(new_n915), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n817), .B1(new_n951), .B2(new_n952), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(KEYINPUT110), .A3(new_n954), .A4(new_n962), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n930), .A2(new_n947), .A3(new_n953), .A4(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n958), .A2(new_n961), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n975), .A3(new_n954), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n971), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g558(.A1(G299), .A2(new_n621), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n587), .B1(new_n615), .B2(new_n620), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT41), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT41), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n622), .A2(new_n587), .ZN(new_n988));
  NAND2_X1  g563(.A1(G299), .A2(new_n621), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n903), .B(new_n630), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT113), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n988), .A2(new_n989), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n993), .A2(KEYINPUT113), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(G288), .B(new_n537), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n721), .A2(G290), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n762), .A2(G305), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n1002), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT42), .Z(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n999), .A2(new_n1001), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n998), .B2(new_n1000), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G868), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n901), .A2(G868), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(G295));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1019), .A3(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(G868), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT114), .B1(new_n1022), .B2(new_n1016), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(G331));
  NAND2_X1  g599(.A1(G301), .A2(G168), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G171), .A2(G286), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n900), .A2(new_n902), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n900), .A2(new_n902), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1027), .B(new_n1029), .C1(new_n986), .C2(new_n990), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1027), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n996), .B1(new_n1031), .B2(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1009), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G37), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1009), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT43), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT41), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n995), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n987), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n988), .A2(new_n989), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(new_n1027), .A3(new_n1029), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1032), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1009), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT43), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1034), .A4(new_n1033), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1035), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT43), .A3(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  MUX2_X1   g627(.A(new_n1048), .B(new_n1052), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g628(.A(new_n752), .B(new_n757), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n845), .A2(G2067), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n916), .A2(new_n847), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n817), .B(G1996), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(G290), .B(new_n764), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1384), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n925), .A2(new_n926), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n489), .A2(G40), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(new_n476), .A3(new_n478), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1063), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1068), .A2(new_n476), .A3(new_n478), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1064), .B1(new_n509), .B2(new_n515), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G305), .A2(G1981), .ZN(new_n1077));
  INV_X1    g652(.A(G1981), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n595), .A2(new_n1078), .A3(new_n601), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(KEYINPUT49), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n545), .A2(G86), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n522), .A2(G48), .ZN(new_n1083));
  AND4_X1   g658(.A1(new_n1078), .A2(new_n1082), .A3(new_n601), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n595), .B2(new_n601), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1086), .A3(new_n1076), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G288), .A2(G1976), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1076), .B1(new_n1089), .B2(new_n1084), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n729), .A2(G1976), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1076), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1093), .B2(KEYINPUT118), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1076), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT119), .B(new_n1091), .C1(new_n729), .C2(G1976), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1976), .B1(new_n591), .B2(new_n593), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(KEYINPUT52), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1097), .B(new_n1087), .C1(new_n1093), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1971), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1069), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT45), .A4(new_n1064), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1074), .A2(KEYINPUT50), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1074), .A2(KEYINPUT50), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(new_n859), .A3(new_n1073), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1104), .A2(new_n1107), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1072), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G303), .A2(G8), .ZN(new_n1115));
  NOR2_X1   g690(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(new_n1116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1090), .B1(new_n1103), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT120), .B1(new_n1123), .B2(new_n1103), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1074), .A2(new_n1066), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1064), .A2(KEYINPUT45), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1073), .B(new_n1126), .C1(G164), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1966), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1108), .A2(new_n1073), .A3(new_n1109), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(G2084), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(G8), .A3(G168), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1125), .B(new_n1133), .C1(new_n1120), .C2(new_n1114), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1087), .B1(new_n1093), .B2(new_n1102), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1096), .B2(new_n1094), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1136), .B(new_n1137), .C1(new_n1120), .C2(new_n1114), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1124), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1131), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1140), .A2(new_n859), .B1(new_n1107), .B2(new_n1104), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1119), .B(new_n1117), .C1(new_n1141), .C2(new_n1072), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1121), .A2(new_n1136), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1125), .B1(new_n1143), .B2(new_n1133), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1122), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G168), .A2(new_n1072), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1132), .B2(G8), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1146), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT51), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(G8), .B(new_n1150), .C1(new_n1132), .C2(G286), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1132), .A2(new_n1146), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1147), .A2(new_n1151), .B1(new_n1132), .B2(new_n1146), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(KEYINPUT126), .A3(new_n1153), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1956), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1131), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(new_n880), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1105), .A2(new_n1106), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n587), .B(KEYINPUT57), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(KEYINPUT122), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1169), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1069), .A2(G2067), .A3(new_n1074), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1131), .B2(new_n806), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n621), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1167), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(G1996), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1106), .A2(new_n1073), .A3(new_n1177), .A4(new_n1126), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT58), .B(G1341), .Z(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1178), .A2(KEYINPUT123), .A3(new_n1180), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n893), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1166), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1168), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1188), .A2(KEYINPUT124), .A3(new_n1167), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n1188), .B2(KEYINPUT124), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n622), .B(new_n1173), .C1(new_n1131), .C2(new_n806), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT60), .B1(new_n1175), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1167), .A2(KEYINPUT61), .B1(new_n1174), .B2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1194), .B(new_n1196), .C1(new_n1185), .C2(KEYINPUT59), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1176), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT53), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1128), .A2(new_n1199), .A3(G2078), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1199), .B1(new_n1107), .B2(G2078), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1131), .A2(new_n793), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(G301), .B(KEYINPUT54), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1204), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1069), .A2(new_n1199), .A3(G2078), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1067), .A2(new_n1207), .A3(new_n1106), .ZN(new_n1208));
  AND4_X1   g783(.A1(new_n1201), .A2(new_n1202), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1143), .A2(new_n1205), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1160), .A2(new_n1198), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1145), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1203), .A2(G171), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1143), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n1215));
  AND3_X1   g790(.A1(new_n1158), .A2(KEYINPUT126), .A3(new_n1153), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT126), .B1(new_n1158), .B2(new_n1153), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1157), .A2(KEYINPUT62), .A3(new_n1159), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1214), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1071), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1070), .A2(new_n764), .A3(new_n762), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT48), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1070), .ZN(new_n1226));
  OAI211_X1 g801(.A(new_n1224), .B(new_n1225), .C1(new_n1061), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1058), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1070), .B1(new_n1229), .B2(new_n915), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1070), .A2(new_n1177), .ZN(new_n1231));
  AND2_X1   g806(.A1(new_n1231), .A2(KEYINPUT46), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1231), .A2(KEYINPUT46), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g809(.A(new_n1234), .B(KEYINPUT47), .Z(new_n1235));
  NAND2_X1  g810(.A1(new_n753), .A2(new_n757), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1057), .B1(new_n1060), .B2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g812(.A(new_n1228), .B(new_n1235), .C1(new_n1070), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1221), .A2(new_n1238), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g814(.A(G319), .B1(new_n662), .B2(new_n663), .ZN(new_n1241));
  NOR2_X1   g815(.A1(G227), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g816(.A1(new_n713), .A2(new_n717), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1243), .B1(new_n1037), .B2(new_n1047), .ZN(new_n1244));
  AOI21_X1  g818(.A(KEYINPUT127), .B1(new_n982), .B2(new_n1244), .ZN(new_n1245));
  AND3_X1   g819(.A1(new_n971), .A2(new_n977), .A3(new_n980), .ZN(new_n1246));
  AOI21_X1  g820(.A(new_n980), .B1(new_n971), .B2(new_n977), .ZN(new_n1247));
  OAI211_X1 g821(.A(KEYINPUT127), .B(new_n1244), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  INV_X1    g822(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g823(.A1(new_n1245), .A2(new_n1249), .ZN(G308));
  OAI21_X1  g824(.A(new_n1244), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1251));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1252));
  NAND2_X1  g826(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n1253), .A2(new_n1248), .ZN(G225));
endmodule


