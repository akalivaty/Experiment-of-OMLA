//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n203), .B1(G155gat), .B2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n205));
  AND2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n202), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n207), .B(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  XOR2_X1   g011(.A(G127gat), .B(G134gat), .Z(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT4), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n217), .ZN(new_n219));
  INV_X1    g018(.A(new_n214), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G225gat), .A2(G233gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(KEYINPUT39), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n210), .B(new_n214), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n225), .B(KEYINPUT39), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G57gat), .B(G85gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT70), .ZN(new_n230));
  XOR2_X1   g029(.A(KEYINPUT69), .B(KEYINPUT0), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G1gat), .B(G29gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(KEYINPUT74), .Z(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT40), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n227), .A2(new_n224), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n222), .B2(new_n224), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n216), .A2(KEYINPUT5), .A3(new_n223), .A4(new_n221), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n243), .A2(new_n235), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n236), .A2(new_n237), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(G183gat), .B(G190gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n249), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n248), .B1(new_n252), .B2(KEYINPUT64), .ZN(new_n253));
  INV_X1    g052(.A(G169gat), .ZN(new_n254));
  INV_X1    g053(.A(G176gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT23), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n253), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  NOR3_X1   g067(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n259), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT67), .B(G197gat), .ZN(new_n278));
  INV_X1    g077(.A(G204gat), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  INV_X1    g080(.A(G211gat), .ZN(new_n282));
  INV_X1    g081(.A(G218gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI22_X1  g083(.A1(new_n280), .A2(new_n281), .B1(KEYINPUT22), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G211gat), .B(G218gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n273), .A2(G226gat), .A3(G233gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n277), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n277), .B2(new_n288), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  OR4_X1    g094(.A1(KEYINPUT30), .A2(new_n290), .A3(new_n291), .A4(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n290), .B2(new_n291), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n289), .A3(new_n294), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n299), .A3(KEYINPUT30), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n274), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n210), .B1(new_n303), .B2(new_n217), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n287), .B1(new_n274), .B2(new_n219), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307));
  OAI211_X1 g106(.A(G228gat), .B(G233gat), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n308), .ZN(new_n310));
  AOI21_X1  g109(.A(G22gat), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(G22gat), .A3(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT31), .B(G50gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n312), .A2(new_n318), .A3(new_n313), .A4(new_n317), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n247), .A2(new_n302), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OR3_X1    g121(.A1(new_n290), .A2(KEYINPUT37), .A3(new_n291), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT75), .B(KEYINPUT38), .Z(new_n324));
  OAI21_X1  g123(.A(KEYINPUT37), .B1(new_n290), .B2(new_n291), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n295), .A4(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n234), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT6), .B1(new_n243), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n244), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n234), .A4(new_n242), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n326), .A2(new_n329), .A3(new_n330), .A4(new_n299), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n323), .A2(new_n295), .A3(new_n325), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n331), .A2(new_n332), .B1(new_n324), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n331), .A2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT77), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n322), .B(new_n338), .C1(new_n334), .C2(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n321), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT73), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n241), .A2(new_n234), .A3(new_n242), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n330), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n301), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n346), .A3(new_n321), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT33), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n273), .A2(new_n220), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n262), .A2(new_n214), .A3(new_n272), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G227gat), .ZN(new_n353));
  INV_X1    g152(.A(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n349), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G15gat), .B(G43gat), .Z(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n350), .A2(new_n351), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n364), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT34), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n352), .B2(new_n356), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n363), .A2(KEYINPUT34), .A3(new_n355), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n365), .B2(new_n366), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT36), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n365), .A2(new_n366), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT66), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n372), .B2(new_n373), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(KEYINPUT66), .A3(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n379), .B2(KEYINPUT36), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n337), .A2(new_n339), .A3(new_n348), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n345), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n377), .A2(new_n340), .A3(new_n382), .A4(new_n378), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT35), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n372), .A2(new_n373), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT35), .B1(new_n329), .B2(new_n330), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n340), .A3(new_n301), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n394));
  NAND2_X1  g193(.A1(G229gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G15gat), .B(G22gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n397), .B2(G1gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G8gat), .ZN(new_n399));
  INV_X1    g198(.A(G1gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(G1gat), .B2(new_n397), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n399), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G43gat), .A2(G50gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G43gat), .A2(G50gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT15), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G29gat), .ZN(new_n410));
  INV_X1    g209(.A(G29gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT80), .B(G36gat), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  OR3_X1    g212(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G36gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n409), .A2(G29gat), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT80), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n408), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n421), .A2(KEYINPUT80), .B1(new_n415), .B2(new_n414), .ZN(new_n424));
  AND2_X1   g223(.A1(KEYINPUT82), .A2(G50gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(KEYINPUT82), .A2(G50gat), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n425), .A2(new_n426), .A3(G43gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT15), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT15), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n431), .A3(new_n405), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n408), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT79), .B(G29gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n434), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n424), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n423), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n404), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n413), .A3(new_n416), .ZN(new_n440));
  OR2_X1    g239(.A1(G43gat), .A2(G50gat), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n430), .B1(new_n441), .B2(new_n405), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n429), .A2(new_n431), .A3(new_n405), .ZN(new_n443));
  INV_X1    g242(.A(new_n426), .ZN(new_n444));
  INV_X1    g243(.A(G43gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(KEYINPUT82), .A2(G50gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n442), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n442), .B1(new_n424), .B2(new_n436), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT17), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n423), .A2(new_n437), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n404), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n451), .A2(new_n404), .A3(KEYINPUT84), .A4(new_n453), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n396), .B(new_n439), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n394), .B1(new_n458), .B2(KEYINPUT18), .ZN(new_n459));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G197gat), .ZN(new_n461));
  XOR2_X1   g260(.A(KEYINPUT11), .B(G169gat), .Z(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT12), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n404), .A2(new_n438), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n404), .A2(new_n438), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n395), .B(KEYINPUT13), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n458), .B2(KEYINPUT18), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n423), .A2(new_n437), .A3(new_n452), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n452), .B1(new_n423), .B2(new_n437), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT84), .B1(new_n475), .B2(new_n404), .ZN(new_n476));
  INV_X1    g275(.A(new_n457), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n395), .B(new_n466), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT18), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n459), .B(new_n465), .C1(new_n472), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n458), .A2(KEYINPUT18), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n468), .A2(new_n470), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n478), .B2(new_n479), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT85), .B1(new_n478), .B2(new_n479), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n464), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G230gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n354), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491));
  INV_X1    g290(.A(G71gat), .ZN(new_n492));
  INV_X1    g291(.A(G78gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G64gat), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(G57gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(G57gat), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n494), .B(KEYINPUT86), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G57gat), .B(G64gat), .Z(new_n502));
  NAND4_X1  g301(.A1(new_n502), .A2(KEYINPUT86), .A3(new_n499), .A4(new_n494), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n501), .A2(KEYINPUT10), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510));
  INV_X1    g309(.A(G85gat), .ZN(new_n511));
  INV_X1    g310(.A(G92gat), .ZN(new_n512));
  AOI22_X1  g311(.A1(KEYINPUT8), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G99gat), .B(G106gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(KEYINPUT8), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n507), .A3(new_n517), .A4(new_n508), .ZN(new_n518));
  INV_X1    g317(.A(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n515), .A2(new_n520), .A3(KEYINPUT90), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT90), .B1(new_n515), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n504), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT95), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n514), .B1(new_n509), .B2(new_n513), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n518), .A2(new_n519), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n515), .A2(new_n520), .A3(KEYINPUT90), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n504), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT10), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n501), .A2(new_n503), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n513), .A2(KEYINPUT93), .A3(new_n507), .A4(new_n508), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n519), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n515), .A2(KEYINPUT94), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n514), .B1(new_n518), .B2(new_n536), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT94), .A3(new_n538), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n535), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n535), .A2(new_n515), .A3(new_n520), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n534), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n490), .B1(new_n533), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n490), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n544), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n548), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n548), .B2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n449), .A2(new_n450), .ZN(new_n558));
  AND2_X1   g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n558), .A2(new_n530), .B1(KEYINPUT41), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n451), .A2(new_n453), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(new_n530), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT91), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n562), .B(new_n564), .Z(new_n565));
  NOR2_X1   g364(.A1(new_n559), .A2(KEYINPUT41), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT89), .ZN(new_n567));
  XOR2_X1   g366(.A(G134gat), .B(G162gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT92), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(new_n565), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n535), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n404), .B1(new_n575), .B2(new_n535), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT88), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT87), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n580), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n574), .A2(new_n588), .ZN(new_n589));
  NOR4_X1   g388(.A1(new_n393), .A2(new_n488), .A3(new_n557), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n344), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n302), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n594), .A2(G8gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT16), .B(G8gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT42), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(KEYINPUT42), .B2(new_n597), .ZN(G1325gat));
  INV_X1    g398(.A(G15gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n590), .A2(new_n600), .A3(new_n385), .ZN(new_n601));
  INV_X1    g400(.A(new_n380), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n590), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n603), .B2(new_n600), .ZN(G1326gat));
  NAND2_X1  g403(.A1(new_n341), .A2(new_n347), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT43), .B(G22gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(G1327gat));
  NOR2_X1   g408(.A1(new_n393), .A2(new_n488), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n574), .A2(new_n557), .A3(new_n588), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR4_X1   g411(.A1(new_n612), .A2(new_n344), .A3(new_n410), .A4(new_n412), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n613), .A2(KEYINPUT45), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(KEYINPUT45), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n388), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n384), .A2(KEYINPUT96), .A3(new_n387), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n381), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n573), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT44), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n574), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n391), .A2(new_n392), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n557), .ZN(new_n626));
  INV_X1    g425(.A(new_n588), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n487), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n344), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n614), .B(new_n615), .C1(new_n435), .C2(new_n630), .ZN(G1328gat));
  NOR3_X1   g430(.A1(new_n612), .A2(G36gat), .A3(new_n301), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(G36gat), .B1(new_n629), .B2(new_n301), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(G1329gat));
  OAI21_X1  g436(.A(G43gat), .B1(new_n629), .B2(new_n380), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT47), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n610), .A2(new_n445), .A3(new_n385), .A4(new_n611), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n638), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(G1330gat));
  NAND2_X1  g442(.A1(new_n444), .A2(new_n446), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n612), .A2(new_n605), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT48), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n644), .B1(new_n629), .B2(new_n340), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR3_X1    g448(.A1(new_n625), .A2(new_n605), .A3(new_n628), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n645), .B1(new_n650), .B2(new_n644), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(KEYINPUT48), .B2(new_n651), .ZN(G1331gat));
  NOR3_X1   g451(.A1(new_n589), .A2(new_n487), .A3(new_n626), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT97), .Z(new_n654));
  AND2_X1   g453(.A1(new_n619), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n591), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g456(.A(new_n301), .B(KEYINPUT98), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT99), .ZN(new_n662));
  NOR2_X1   g461(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(G1333gat));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n380), .A2(new_n492), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n655), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n655), .B2(new_n666), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n655), .A2(new_n385), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n667), .A2(new_n668), .B1(G71gat), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n606), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT101), .B(G78gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1335gat));
  NOR2_X1   g473(.A1(new_n487), .A2(new_n588), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n625), .A2(new_n626), .A3(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(new_n591), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n619), .A2(new_n573), .A3(new_n675), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT51), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n591), .A2(new_n511), .A3(new_n557), .ZN(new_n683));
  OAI22_X1  g482(.A1(new_n678), .A2(new_n511), .B1(new_n682), .B2(new_n683), .ZN(G1336gat));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n658), .A2(new_n512), .A3(new_n557), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT102), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n676), .A2(new_n626), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n622), .A2(new_n624), .A3(new_n658), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G92gat), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT52), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n622), .A2(new_n624), .A3(new_n302), .A4(new_n689), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G92gat), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n688), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n685), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n688), .A2(new_n696), .ZN(new_n699));
  OAI211_X1 g498(.A(KEYINPUT103), .B(new_n693), .C1(new_n699), .C2(new_n692), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1337gat));
  INV_X1    g500(.A(G99gat), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n681), .A2(new_n702), .A3(new_n385), .A4(new_n557), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n677), .A2(new_n602), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n702), .ZN(G1338gat));
  INV_X1    g504(.A(G106gat), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n677), .B2(new_n606), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n340), .A2(G106gat), .A3(new_n626), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n681), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT53), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n340), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n622), .A2(new_n624), .A3(new_n711), .A4(new_n689), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n706), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n392), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT78), .B1(new_n381), .B2(new_n388), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n717), .A2(new_n623), .B1(new_n621), .B2(new_n620), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n718), .A2(KEYINPUT105), .A3(new_n711), .A4(new_n689), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT104), .B(KEYINPUT53), .Z(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n681), .B2(new_n708), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n720), .A2(KEYINPUT106), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT106), .B1(new_n720), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n710), .B1(new_n723), .B2(new_n724), .ZN(G1339gat));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n501), .A2(KEYINPUT10), .A3(new_n503), .ZN(new_n727));
  AOI211_X1 g526(.A(KEYINPUT95), .B(new_n727), .C1(new_n528), .C2(new_n529), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n531), .B1(new_n530), .B2(new_n504), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n501), .A2(new_n503), .ZN(new_n731));
  INV_X1    g530(.A(new_n543), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n542), .A2(new_n538), .B1(new_n515), .B2(KEYINPUT94), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT10), .B1(new_n734), .B2(new_n545), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n549), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n533), .A2(new_n547), .A3(new_n490), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(KEYINPUT54), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT54), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n553), .B1(new_n548), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n740), .A3(KEYINPUT55), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n555), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT55), .B1(new_n738), .B2(new_n740), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n487), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n484), .A2(new_n464), .A3(new_n482), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n456), .A2(new_n457), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n395), .B1(new_n750), .B2(new_n466), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n463), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n746), .A2(new_n557), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n573), .B1(new_n745), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n573), .A2(new_n744), .A3(new_n746), .A4(new_n752), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n726), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n746), .A2(new_n557), .A3(new_n752), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n487), .B2(new_n744), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT108), .B(new_n755), .C1(new_n759), .C2(new_n573), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n627), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n488), .A2(new_n574), .A3(new_n626), .A4(new_n588), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n658), .A2(new_n344), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(new_n605), .A3(new_n385), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(G113gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n769), .A2(new_n770), .A3(new_n488), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n767), .A2(new_n591), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n379), .A2(new_n711), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(new_n659), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n774), .A2(new_n488), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n771), .B1(new_n775), .B2(new_n770), .ZN(G1340gat));
  OAI21_X1  g575(.A(G120gat), .B1(new_n769), .B2(new_n626), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n626), .A2(G120gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT110), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n774), .B2(new_n779), .ZN(G1341gat));
  INV_X1    g579(.A(G127gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n769), .A2(new_n781), .A3(new_n627), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n774), .A2(KEYINPUT111), .A3(new_n627), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(G127gat), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT111), .B1(new_n774), .B2(new_n627), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(G1342gat));
  NAND2_X1  g585(.A1(new_n301), .A2(new_n573), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(G134gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT56), .ZN(new_n790));
  OAI21_X1  g589(.A(G134gat), .B1(new_n769), .B2(new_n574), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(KEYINPUT56), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(G1343gat));
  NOR2_X1   g592(.A1(new_n602), .A2(new_n340), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n658), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n488), .A2(G141gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n767), .A2(new_n800), .A3(new_n711), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n380), .A2(new_n768), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n380), .A2(new_n768), .A3(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n738), .B2(new_n740), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n742), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n758), .B1(new_n487), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n755), .B1(new_n810), .B2(new_n573), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n627), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n762), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n812), .A2(KEYINPUT114), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n606), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n806), .B1(KEYINPUT57), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G141gat), .B1(new_n818), .B2(new_n488), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT58), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT58), .B1(new_n797), .B2(new_n798), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT117), .A3(new_n819), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT117), .B1(new_n824), .B2(new_n819), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G1344gat));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828));
  INV_X1    g627(.A(G148gat), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n340), .A2(new_n800), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n764), .A2(new_n766), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n764), .A2(KEYINPUT118), .A3(new_n766), .A4(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n812), .A2(new_n762), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT119), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n605), .B1(new_n835), .B2(KEYINPUT119), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n800), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n806), .A2(new_n626), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n828), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n841), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n831), .A2(new_n832), .B1(new_n838), .B2(new_n800), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n834), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n847), .C2(new_n829), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n818), .A2(new_n626), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n843), .A2(G148gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n797), .A2(new_n829), .A3(new_n557), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(KEYINPUT121), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n852), .B1(new_n844), .B2(new_n848), .ZN(new_n858));
  INV_X1    g657(.A(new_n855), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(G1345gat));
  INV_X1    g660(.A(G155gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n797), .A2(new_n862), .A3(new_n588), .ZN(new_n863));
  OAI21_X1  g662(.A(G155gat), .B1(new_n818), .B2(new_n627), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n818), .B2(new_n574), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n787), .A2(G162gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n796), .B2(new_n867), .ZN(G1347gat));
  AND2_X1   g667(.A1(new_n767), .A2(new_n344), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n659), .A2(new_n379), .A3(new_n711), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(G169gat), .A3(new_n488), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n302), .A2(new_n344), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n372), .A3(new_n373), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT123), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n767), .A2(new_n605), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n488), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n878), .ZN(G1348gat));
  OAI21_X1  g678(.A(G176gat), .B1(new_n877), .B2(new_n626), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n557), .A2(new_n255), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n871), .B2(new_n881), .ZN(G1349gat));
  NOR2_X1   g681(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n883));
  OR3_X1    g682(.A1(new_n877), .A2(KEYINPUT124), .A3(new_n627), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n877), .B2(new_n627), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(G183gat), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n263), .A3(new_n588), .A4(new_n870), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n877), .B2(new_n574), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT61), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n573), .A2(new_n264), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n871), .B2(new_n893), .ZN(G1351gat));
  NAND2_X1  g693(.A1(new_n794), .A2(new_n658), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT126), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n869), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G197gat), .B1(new_n898), .B2(new_n487), .ZN(new_n899));
  INV_X1    g698(.A(new_n840), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n602), .A2(new_n874), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n487), .A2(G197gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(G1352gat));
  NOR3_X1   g704(.A1(new_n897), .A2(G204gat), .A3(new_n626), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT62), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n900), .A2(new_n626), .A3(new_n902), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n279), .B2(new_n908), .ZN(G1353gat));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n282), .A3(new_n588), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n903), .A2(new_n588), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n282), .B1(KEYINPUT127), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n912), .A2(new_n915), .B1(new_n911), .B2(KEYINPUT63), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n913), .B2(new_n916), .ZN(G1354gat));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n283), .A3(new_n573), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n900), .A2(new_n574), .A3(new_n902), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n283), .ZN(G1355gat));
endmodule


