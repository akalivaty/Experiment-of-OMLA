//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(G50gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(G43gat), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n205), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT82), .B(G43gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT14), .B(G29gat), .Z(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G36gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n208), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n208), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G8gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n226), .B(G8gat), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT84), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT84), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n214), .A2(new_n218), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n234), .B(new_n220), .C1(new_n235), .C2(new_n208), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT17), .B1(new_n219), .B2(new_n221), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n203), .B(new_n228), .C1(new_n233), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n202), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G197gat), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT11), .B(G169gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n203), .B(KEYINPUT13), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n220), .B1(new_n235), .B2(new_n208), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n229), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n251), .B2(new_n228), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n239), .B2(new_n240), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n236), .A2(new_n237), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n232), .A3(new_n230), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n255), .A2(KEYINPUT18), .A3(new_n203), .A4(new_n228), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n253), .B(new_n256), .C1(new_n241), .C2(new_n246), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G183gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT27), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT27), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT27), .B(G183gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT28), .A3(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT26), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n265), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n269), .A2(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n288));
  OR3_X1    g087(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n276), .B2(KEYINPUT24), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND4_X1   g093(.A1(KEYINPUT25), .A2(new_n288), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n287), .B2(KEYINPUT24), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT25), .B1(new_n296), .B2(new_n291), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n284), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT64), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT65), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(KEYINPUT1), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(G134gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n304), .B2(KEYINPUT1), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G134gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(G120gat), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n316), .B(new_n303), .C1(new_n306), .C2(new_n308), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n310), .A2(new_n317), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n288), .A2(new_n291), .A3(new_n294), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n291), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n325), .A3(new_n284), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n319), .A2(new_n326), .A3(G227gat), .A4(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT33), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n264), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(KEYINPUT32), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(KEYINPUT66), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT33), .B1(new_n264), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n335), .B2(new_n264), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n326), .ZN(new_n341));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n333), .A2(new_n340), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n344), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n329), .A2(new_n330), .B1(KEYINPUT32), .B2(new_n327), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n329), .B2(KEYINPUT66), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G22gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT2), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G155gat), .B(G162gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G141gat), .B(G148gat), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n354), .A2(KEYINPUT2), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G148gat), .ZN(new_n363));
  INV_X1    g162(.A(G148gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G141gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n355), .B(new_n366), .C1(new_n369), .C2(new_n356), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n361), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n361), .A2(new_n370), .A3(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G197gat), .ZN(new_n376));
  INV_X1    g175(.A(G204gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  NAND2_X1  g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n378), .A2(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n380), .ZN(new_n385));
  NOR2_X1   g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386));
  AND2_X1   g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n381), .ZN(new_n389));
  NOR2_X1   g188(.A1(G211gat), .A2(G218gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT3), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n375), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n371), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT74), .B(KEYINPUT3), .C1(new_n361), .C2(new_n370), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n393), .B(KEYINPUT69), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(new_n405), .B2(KEYINPUT79), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n353), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n382), .B2(new_n383), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT77), .B1(new_n388), .B2(new_n391), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n388), .A2(KEYINPUT78), .A3(new_n391), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n382), .A2(new_n414), .A3(new_n383), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT3), .B1(new_n416), .B2(new_n397), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n353), .B1(new_n417), .B2(new_n371), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n404), .B2(new_n402), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n352), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n397), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n371), .A2(new_n399), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT74), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n371), .A2(new_n398), .A3(new_n399), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT79), .B1(new_n425), .B2(new_n403), .ZN(new_n426));
  INV_X1    g225(.A(new_n396), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n408), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n353), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n419), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(G22gat), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT31), .B(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n420), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n420), .B2(new_n432), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n351), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G8gat), .B(G36gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  AND2_X1   g240(.A1(new_n441), .A2(KEYINPUT30), .ZN(new_n442));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n298), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n325), .A2(KEYINPUT70), .A3(new_n284), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n298), .A2(new_n394), .A3(new_n443), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n447), .A2(new_n449), .A3(new_n404), .ZN(new_n450));
  INV_X1    g249(.A(new_n443), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n421), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n325), .A2(new_n284), .A3(new_n451), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n403), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n442), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n404), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n298), .A2(new_n444), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT70), .B1(new_n325), .B2(new_n284), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n451), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n403), .A3(new_n448), .ZN(new_n462));
  INV_X1    g261(.A(new_n441), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n458), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n456), .B(new_n464), .C1(new_n465), .C2(KEYINPUT30), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT0), .ZN(new_n469));
  XNOR2_X1  g268(.A(G57gat), .B(G85gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n471), .A2(KEYINPUT6), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n361), .A2(new_n370), .A3(KEYINPUT73), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT73), .B1(new_n361), .B2(new_n370), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n318), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI221_X4 g277(.A(KEYINPUT75), .B1(new_n361), .B2(new_n370), .C1(new_n310), .C2(new_n317), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT75), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n318), .B2(new_n371), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT76), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n318), .A2(new_n371), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT75), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n318), .A2(new_n480), .A3(new_n371), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n373), .A2(KEYINPUT3), .A3(new_n374), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(new_n320), .C1(new_n400), .C2(new_n401), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n318), .A2(KEYINPUT4), .A3(new_n371), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n489), .A2(new_n491), .A3(new_n483), .A4(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n373), .A2(new_n317), .A3(new_n310), .A4(new_n374), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n486), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT76), .ZN(new_n496));
  INV_X1    g295(.A(new_n483), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n484), .A2(KEYINPUT5), .A3(new_n493), .A4(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n491), .A2(new_n483), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n487), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT4), .B1(new_n479), .B2(new_n481), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AOI211_X1 g303(.A(new_n474), .B(new_n475), .C1(new_n499), .C2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n499), .A2(new_n473), .A3(new_n504), .A4(new_n472), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT81), .B(new_n467), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT35), .B1(new_n438), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n435), .ZN(new_n510));
  AOI21_X1  g309(.A(G22gat), .B1(new_n430), .B2(new_n431), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n352), .B(new_n419), .C1(new_n428), .C2(new_n429), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n420), .A2(new_n432), .A3(new_n435), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n513), .A2(new_n514), .B1(new_n346), .B2(new_n350), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n504), .ZN(new_n517));
  INV_X1    g316(.A(new_n474), .ZN(new_n518));
  INV_X1    g317(.A(new_n475), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n466), .B1(new_n520), .B2(new_n506), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n515), .A2(KEYINPUT81), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n509), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n458), .A2(KEYINPUT37), .A3(new_n462), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n450), .A2(new_n455), .A3(new_n441), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n463), .A2(KEYINPUT37), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT38), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n453), .A2(new_n454), .A3(new_n403), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n530), .A2(KEYINPUT37), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n404), .B1(new_n447), .B2(new_n449), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT38), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n464), .A2(new_n526), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n465), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n529), .A2(new_n535), .A3(new_n520), .A4(new_n506), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n514), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT40), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n503), .A2(new_n491), .A3(new_n502), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n497), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n486), .A2(new_n483), .A3(new_n488), .A4(new_n494), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT39), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT80), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(KEYINPUT80), .A3(KEYINPUT39), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(new_n547), .A3(new_n497), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n471), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n538), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n517), .A2(new_n472), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(KEYINPUT40), .A3(new_n471), .A4(new_n548), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n466), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n436), .A2(new_n437), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n467), .B1(new_n505), .B2(new_n507), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n351), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT68), .B(KEYINPUT36), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n346), .A2(new_n350), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n261), .B1(new_n523), .B2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G57gat), .B(G64gat), .Z(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(KEYINPUT87), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT86), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n229), .B1(new_n575), .B2(new_n576), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT88), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n581), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT89), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT91), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n600), .A2(new_n603), .A3(new_n604), .A4(new_n596), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n599), .B(new_n605), .C1(new_n606), .C2(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n608), .B1(new_n601), .B2(new_n602), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G99gat), .B(G106gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT92), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n611), .B(KEYINPUT92), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n607), .A3(new_n609), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(KEYINPUT93), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT93), .B1(new_n613), .B2(new_n615), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n254), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n610), .A2(new_n612), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n614), .B1(new_n607), .B2(new_n609), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n616), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT94), .B1(new_n626), .B2(new_n238), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n626), .A2(new_n222), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT95), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n619), .B2(new_n250), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n627), .B2(new_n621), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT96), .B1(new_n636), .B2(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n628), .A2(new_n631), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n629), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n595), .B1(new_n633), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n632), .B(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n644), .A2(new_n637), .A3(new_n640), .A4(new_n594), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n573), .B(new_n574), .Z(new_n648));
  NOR2_X1   g447(.A1(new_n623), .A2(new_n624), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n610), .A2(KEYINPUT97), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  OAI22_X1  g451(.A1(new_n575), .A2(new_n650), .B1(new_n623), .B2(new_n624), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  AOI211_X1 g454(.A(new_n655), .B(new_n575), .C1(new_n625), .C2(new_n616), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n647), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  INV_X1    g457(.A(new_n647), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n657), .A2(new_n660), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n657), .B2(new_n660), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n565), .A2(new_n588), .A3(new_n646), .A4(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(KEYINPUT99), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(KEYINPUT99), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n505), .A2(new_n507), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  NAND4_X1  g476(.A1(new_n673), .A2(KEYINPUT42), .A3(new_n466), .A4(new_n677), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n672), .A2(KEYINPUT100), .A3(new_n467), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT100), .B1(new_n672), .B2(new_n467), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(G8gat), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n677), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n678), .B(new_n681), .C1(new_n683), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n672), .B2(new_n563), .ZN(new_n685));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n351), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n672), .B2(new_n687), .ZN(G1326gat));
  OR3_X1    g487(.A1(new_n672), .A2(KEYINPUT101), .A3(new_n537), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT101), .B1(new_n672), .B2(new_n537), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NOR3_X1   g492(.A1(new_n438), .A2(new_n508), .A3(KEYINPUT35), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT81), .ZN(new_n695));
  AOI211_X1 g494(.A(new_n695), .B(new_n466), .C1(new_n520), .C2(new_n506), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n516), .B1(new_n696), .B2(new_n515), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n564), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n642), .A2(new_n645), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n537), .B2(new_n521), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT104), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n555), .A4(new_n563), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n523), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n642), .A2(new_n645), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n702), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  AOI211_X1 g510(.A(KEYINPUT105), .B(new_n709), .C1(new_n706), .C2(new_n523), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n701), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n668), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n588), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n261), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT103), .Z(new_n718));
  AND2_X1   g517(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n674), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n700), .A2(new_n261), .A3(new_n716), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n215), .A3(new_n674), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(G1328gat));
  INV_X1    g526(.A(G36gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(new_n728), .A3(new_n466), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n720), .B2(new_n467), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(G1329gat));
  OR3_X1    g534(.A1(new_n720), .A2(new_n563), .A3(new_n212), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n351), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n212), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1330gat));
  OAI21_X1  g542(.A(G50gat), .B1(new_n720), .B2(new_n537), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n716), .A2(G50gat), .A3(new_n537), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n565), .A2(new_n699), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1331gat));
  INV_X1    g548(.A(new_n588), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n699), .A2(new_n260), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n714), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n707), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n674), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n467), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g560(.A(G64gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n755), .A2(new_n763), .A3(new_n759), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n758), .A2(new_n761), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n761), .A2(new_n764), .B1(new_n758), .B2(new_n762), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(G1333gat));
  NAND2_X1  g566(.A1(new_n755), .A2(new_n351), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n568), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n563), .A2(new_n568), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n755), .B2(new_n771), .ZN(new_n772));
  AND4_X1   g571(.A1(new_n770), .A2(new_n754), .A3(new_n707), .A4(new_n771), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n769), .B(new_n775), .C1(new_n772), .C2(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n755), .A2(new_n556), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g580(.A1(new_n750), .A2(new_n261), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n646), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n707), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n668), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n601), .A3(new_n674), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n782), .A2(new_n668), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n713), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G85gat), .B1(new_n794), .B2(new_n721), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1336gat));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n713), .A2(new_n466), .A3(new_n793), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n668), .A2(G92gat), .A3(new_n467), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n797), .B(new_n799), .C1(new_n790), .C2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  INV_X1    g602(.A(new_n785), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n799), .A2(new_n803), .B1(new_n804), .B2(new_n800), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n798), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n806));
  AOI211_X1 g605(.A(KEYINPUT114), .B(new_n797), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n799), .A2(new_n803), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n800), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(KEYINPUT52), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n802), .B1(new_n807), .B2(new_n812), .ZN(G1337gat));
  INV_X1    g612(.A(G99gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n791), .A2(new_n814), .A3(new_n351), .ZN(new_n815));
  OAI21_X1  g614(.A(G99gat), .B1(new_n794), .B2(new_n563), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n794), .B2(new_n537), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n537), .A2(G106gat), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n786), .A2(new_n714), .A3(new_n789), .A4(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(KEYINPUT116), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(KEYINPUT116), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n818), .B(new_n819), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n804), .A2(new_n714), .A3(new_n820), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n818), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n647), .C1(new_n654), .C2(new_n656), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n664), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n648), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n659), .B(new_n834), .C1(new_n658), .C2(KEYINPUT10), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n836), .A3(KEYINPUT55), .ZN(new_n837));
  INV_X1    g636(.A(new_n666), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n228), .B1(new_n233), .B2(new_n238), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(G229gat), .A3(G233gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n251), .A2(new_n228), .A3(new_n249), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT118), .Z(new_n845));
  NAND4_X1  g644(.A1(new_n840), .A2(KEYINPUT117), .A3(G229gat), .A4(G233gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n257), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n847), .A2(new_n245), .B1(new_n848), .B2(new_n246), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT55), .B1(new_n833), .B2(new_n836), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n839), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n646), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n851), .A2(new_n260), .A3(new_n838), .A4(new_n837), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n714), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n854), .A2(new_n855), .B1(new_n642), .B2(new_n645), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n750), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n646), .A2(new_n261), .A3(new_n588), .A4(new_n668), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n721), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n438), .A2(new_n466), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n260), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n515), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n721), .A2(new_n466), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n261), .A2(new_n312), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(G1340gat));
  AOI21_X1  g669(.A(G120gat), .B1(new_n862), .B2(new_n714), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n668), .A2(new_n314), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n868), .B2(new_n872), .ZN(G1341gat));
  INV_X1    g672(.A(new_n868), .ZN(new_n874));
  OAI21_X1  g673(.A(G127gat), .B1(new_n874), .B2(new_n750), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n750), .A2(G127gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n861), .B2(new_n876), .ZN(G1342gat));
  NOR3_X1   g676(.A1(new_n861), .A2(G134gat), .A3(new_n646), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n874), .B2(new_n646), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  NAND2_X1  g682(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n884));
  INV_X1    g683(.A(new_n563), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n466), .A3(new_n537), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n859), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n261), .A2(G141gat), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n884), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n867), .A2(new_n885), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT119), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n847), .A2(new_n245), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n848), .A2(new_n246), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n850), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(new_n642), .A3(new_n645), .A4(new_n839), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n668), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n850), .B(new_n899), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n260), .A2(new_n838), .A3(new_n837), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n897), .B1(new_n902), .B2(new_n699), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n903), .A2(new_n750), .B1(new_n668), .B2(new_n751), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n537), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n864), .B2(new_n556), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n260), .B(new_n892), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n890), .B1(new_n908), .B2(G141gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(G1344gat));
  OAI21_X1  g710(.A(KEYINPUT59), .B1(new_n887), .B2(new_n668), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n364), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n906), .A2(new_n907), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n892), .A2(new_n714), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT59), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n905), .B1(new_n904), .B2(new_n537), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n556), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n920));
  OAI221_X1 g719(.A(new_n913), .B1(new_n914), .B2(new_n916), .C1(new_n919), .C2(new_n920), .ZN(G1345gat));
  INV_X1    g720(.A(new_n892), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n588), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G155gat), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n750), .A2(G155gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n887), .B2(new_n926), .ZN(G1346gat));
  INV_X1    g726(.A(G162gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n646), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n859), .A2(new_n699), .A3(new_n886), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n923), .A2(new_n929), .B1(new_n928), .B2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n674), .A2(new_n467), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n864), .A2(new_n515), .A3(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(new_n277), .A3(new_n261), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n864), .A2(new_n721), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n864), .A2(new_n937), .A3(new_n721), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n515), .A2(new_n466), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT123), .Z(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n260), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n934), .B1(new_n942), .B2(new_n277), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n933), .B2(new_n668), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n714), .A2(new_n278), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n933), .B2(new_n750), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n588), .A2(new_n273), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g750(.A1(new_n939), .A2(new_n269), .A3(new_n699), .A4(new_n941), .ZN(new_n952));
  OAI21_X1  g751(.A(G190gat), .B1(new_n933), .B2(new_n646), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n952), .B(KEYINPUT124), .C1(new_n955), .C2(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1351gat));
  NOR3_X1   g760(.A1(new_n885), .A2(new_n467), .A3(new_n537), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n939), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n260), .ZN(new_n964));
  INV_X1    g763(.A(new_n932), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n885), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n967), .B1(new_n917), .B2(new_n918), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n261), .A2(new_n376), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  AOI21_X1  g769(.A(new_n377), .B1(new_n968), .B2(new_n714), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n668), .A2(G204gat), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n939), .A2(new_n972), .A3(new_n962), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n937), .B1(new_n864), .B2(new_n721), .ZN(new_n975));
  AOI211_X1 g774(.A(KEYINPUT122), .B(new_n674), .C1(new_n857), .C2(new_n858), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n962), .B(new_n973), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n971), .B1(new_n979), .B2(KEYINPUT62), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(KEYINPUT126), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(KEYINPUT126), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(G1353gat));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n903), .A2(new_n750), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n537), .B1(new_n987), .B2(new_n858), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n918), .B1(new_n988), .B2(KEYINPUT57), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n588), .A4(new_n966), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT127), .B1(new_n968), .B2(new_n588), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n989), .A2(new_n588), .A3(new_n966), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n990), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(G211gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n963), .A2(new_n999), .A3(new_n588), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1354gat));
  INV_X1    g800(.A(G218gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n963), .A2(new_n1002), .A3(new_n699), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n968), .A2(new_n699), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n1002), .B2(new_n1004), .ZN(G1355gat));
endmodule


