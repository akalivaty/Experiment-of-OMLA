//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT68), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G107), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n204), .C2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n205), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n204), .A2(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n189), .A2(new_n217), .A3(G143), .A4(new_n190), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT64), .A2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT64), .A2(G146), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n219), .A2(new_n220), .A3(new_n192), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT65), .B1(new_n188), .B2(G143), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(new_n223), .B2(new_n226), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n200), .B(new_n216), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT79), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n194), .A2(KEYINPUT79), .A3(KEYINPUT1), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n232), .A2(G128), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(new_n223), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n219), .A2(new_n220), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n222), .B1(new_n236), .B2(G143), .ZN(new_n237));
  INV_X1    g051(.A(new_n218), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n226), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT67), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n235), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n229), .B1(new_n242), .B2(new_n216), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT11), .B1(new_n244), .B2(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT66), .A2(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT66), .A2(G137), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT11), .A2(G134), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n247), .B2(new_n251), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n243), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT12), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n243), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n211), .A2(new_n208), .A3(new_n203), .A4(new_n205), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G101), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(new_n222), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n196), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n266), .B2(new_n218), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n193), .B2(new_n194), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n261), .A2(new_n272), .A3(G101), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n261), .A2(KEYINPUT78), .A3(new_n272), .A4(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n200), .B1(new_n227), .B2(new_n228), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT10), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n216), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n271), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n242), .B2(new_n216), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n255), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n258), .A2(new_n260), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G110), .B(G140), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G227), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n285), .B(new_n287), .Z(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n255), .B1(new_n281), .B2(new_n282), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n288), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n283), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT80), .A3(G469), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n289), .B2(new_n293), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n278), .A2(new_n280), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n271), .A2(new_n277), .ZN(new_n303));
  AND4_X1   g117(.A1(new_n255), .A2(new_n282), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n288), .B1(new_n304), .B2(new_n290), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n258), .A2(new_n260), .A3(new_n283), .A4(new_n292), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n300), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n297), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G221), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n312), .B2(new_n295), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G210), .B1(G237), .B2(G902), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n316), .B(KEYINPUT85), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G125), .B1(new_n267), .B2(new_n269), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n221), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G128), .A3(new_n197), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n240), .A2(new_n241), .B1(new_n195), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G224), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G953), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT7), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT83), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT8), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n212), .A2(new_n215), .ZN(new_n336));
  INV_X1    g150(.A(G116), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT70), .B1(new_n337), .B2(G119), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n339));
  INV_X1    g153(.A(G119), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT2), .A2(G113), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT2), .ZN(new_n347));
  INV_X1    g161(.A(G113), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(G116), .ZN(new_n353));
  OAI21_X1  g167(.A(G113), .B1(new_n353), .B2(KEYINPUT5), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n338), .A2(new_n341), .A3(KEYINPUT5), .A4(new_n342), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n335), .B1(new_n336), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n354), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n360), .B2(new_n356), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n216), .B1(new_n362), .B2(new_n352), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n358), .A2(new_n216), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n351), .B(new_n343), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(new_n262), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n368), .B2(new_n277), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n364), .B1(new_n369), .B2(new_n334), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n327), .A2(new_n332), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n319), .B1(new_n278), .B2(G125), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n331), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n333), .A2(new_n370), .A3(new_n371), .A4(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n295), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n372), .B(new_n329), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n369), .B2(new_n334), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n334), .B(KEYINPUT81), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n369), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n369), .A2(new_n379), .A3(new_n382), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n376), .B1(new_n375), .B2(new_n295), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n318), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n375), .A2(new_n295), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT84), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(new_n317), .A3(new_n386), .A4(new_n377), .ZN(new_n392));
  OAI21_X1  g206(.A(G214), .B1(G237), .B2(G902), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  NOR2_X1   g210(.A1(G237), .A2(G953), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G214), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n192), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(G143), .A3(G214), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT18), .A3(G131), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n401), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT88), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(KEYINPUT89), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G125), .B(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n236), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n188), .B2(new_n413), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT87), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n404), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n418));
  OR3_X1    g232(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n188), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(G146), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n401), .A2(KEYINPUT17), .A3(G131), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n401), .B(G131), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n424), .B(new_n425), .C1(KEYINPUT17), .C2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n204), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n417), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n413), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT19), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n426), .B(new_n422), .C1(new_n191), .C2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n429), .B1(new_n417), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n395), .B(new_n396), .C1(new_n431), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT91), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n417), .A2(new_n435), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n430), .B1(new_n439), .B2(new_n429), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n395), .A4(new_n396), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n396), .B1(new_n431), .B2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT20), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n429), .B1(new_n417), .B2(new_n427), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n295), .B1(new_n431), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT92), .B(new_n295), .C1(new_n431), .C2(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(G475), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G478), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n192), .A2(G128), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT13), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n192), .B2(G128), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n225), .A2(KEYINPUT93), .A3(G143), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n459), .B1(new_n465), .B2(KEYINPUT94), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(KEYINPUT94), .B2(new_n465), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G134), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n457), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G134), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n337), .A2(G122), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G107), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n202), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n337), .A2(KEYINPUT14), .A3(G122), .ZN(new_n479));
  OAI211_X1 g293(.A(G107), .B(new_n479), .C1(new_n474), .C2(KEYINPUT14), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT95), .Z(new_n481));
  XNOR2_X1  g295(.A(new_n469), .B(G134), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G217), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n311), .A2(new_n485), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n483), .A3(new_n486), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n456), .B1(new_n490), .B2(new_n295), .ZN(new_n491));
  AOI211_X1 g305(.A(G902), .B(new_n455), .C1(new_n488), .C2(new_n489), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n286), .A2(G952), .ZN(new_n495));
  INV_X1    g309(.A(G234), .ZN(new_n496));
  INV_X1    g310(.A(G237), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n295), .B(new_n286), .C1(G234), .C2(G237), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(G898), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n453), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n315), .A2(new_n394), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(G472), .A2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n256), .B2(new_n270), .ZN(new_n511));
  INV_X1    g325(.A(new_n253), .ZN(new_n512));
  AOI21_X1  g326(.A(G134), .B1(new_n248), .B2(new_n249), .ZN(new_n513));
  INV_X1    g327(.A(new_n246), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n511), .B1(new_n325), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n344), .B(new_n351), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n255), .A2(new_n267), .A3(new_n269), .ZN(new_n519));
  INV_X1    g333(.A(new_n516), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n278), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n517), .B(new_n518), .C1(new_n521), .C2(KEYINPUT30), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n397), .A2(G210), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n523), .B(KEYINPUT27), .Z(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n521), .B2(new_n366), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n528), .B2(KEYINPUT31), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  AOI211_X1 g347(.A(KEYINPUT71), .B(new_n533), .C1(new_n522), .C2(new_n527), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n526), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT28), .B1(new_n521), .B2(new_n366), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT28), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n240), .A2(new_n241), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n516), .B1(new_n539), .B2(new_n200), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n518), .B1(new_n540), .B2(new_n519), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n278), .A2(new_n520), .ZN(new_n542));
  INV_X1    g356(.A(new_n519), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n366), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n538), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n537), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n540), .A2(new_n518), .A3(new_n519), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n366), .B1(new_n542), .B2(new_n543), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT28), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n536), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n509), .B1(new_n535), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n545), .A2(new_n537), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n526), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n547), .A2(new_n536), .A3(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n522), .A2(new_n544), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n526), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n556), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n558), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT75), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n509), .C1(new_n535), .C2(new_n552), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n554), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n506), .B1(new_n535), .B2(new_n552), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT74), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n570), .B(new_n506), .C1(new_n535), .C2(new_n552), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n508), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(new_n340), .B2(G128), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n576), .C1(G119), .C2(new_n225), .ZN(new_n577));
  XNOR2_X1  g391(.A(G119), .B(G128), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT24), .B(G110), .Z(new_n579));
  AOI22_X1  g393(.A1(new_n577), .A2(G110), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n423), .A2(new_n580), .ZN(new_n581));
  OAI22_X1  g395(.A1(new_n577), .A2(G110), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n422), .A3(new_n414), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT22), .B(G137), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n310), .A2(new_n496), .A3(G953), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n581), .A2(new_n583), .A3(new_n587), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT25), .B1(new_n591), .B2(new_n295), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(KEYINPUT25), .A3(new_n295), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n485), .B1(G234), .B2(new_n295), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT76), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n591), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n596), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n505), .A2(new_n573), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT96), .B(G101), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  OAI21_X1  g422(.A(new_n295), .B1(new_n535), .B2(new_n552), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n569), .A2(new_n571), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n490), .A2(new_n454), .A3(new_n295), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n454), .B2(new_n295), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n490), .A2(KEYINPUT33), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n488), .A2(new_n489), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n452), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n394), .A2(KEYINPUT98), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n389), .A2(new_n392), .A3(new_n625), .A4(new_n393), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n502), .B(new_n623), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n605), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n315), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n615), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n444), .A2(new_n437), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n444), .A2(KEYINPUT100), .A3(new_n437), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(new_n494), .A3(new_n451), .A4(new_n637), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n502), .B(new_n638), .C1(new_n624), .C2(new_n626), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n615), .A2(new_n639), .A3(new_n629), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n584), .B(new_n643), .Z(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n603), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n595), .B2(new_n599), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n615), .A2(new_n505), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n499), .B1(new_n500), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n638), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n569), .A2(new_n508), .A3(new_n571), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n554), .A2(new_n564), .A3(new_n566), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n647), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n309), .A2(new_n314), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n624), .A2(new_n626), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n225), .ZN(G30));
  NAND2_X1  g476(.A1(new_n389), .A2(new_n392), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n453), .A2(new_n493), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n393), .A2(new_n668), .A3(new_n646), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n652), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n658), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n526), .B1(new_n522), .B2(new_n544), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n541), .A2(new_n526), .A3(new_n544), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n295), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT102), .Z(new_n679));
  AND3_X1   g493(.A1(new_n554), .A2(new_n566), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n572), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n670), .A2(new_n673), .A3(new_n674), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NOR3_X1   g497(.A1(new_n623), .A2(new_n646), .A3(new_n652), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n655), .B2(new_n656), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT103), .B1(new_n685), .B2(new_n660), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n315), .B1(new_n624), .B2(new_n626), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n573), .A4(new_n684), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  OR2_X1    g505(.A1(new_n307), .A2(new_n300), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(KEYINPUT104), .A3(new_n308), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n307), .A2(KEYINPUT104), .A3(new_n300), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n313), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n627), .A2(new_n573), .A3(new_n605), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT105), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n697), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n639), .A2(new_n573), .A3(new_n605), .A4(new_n696), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT106), .B(G116), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G18));
  NOR2_X1   g517(.A1(new_n307), .A2(new_n300), .ZN(new_n704));
  AOI211_X1 g518(.A(G469), .B(G902), .C1(new_n305), .C2(new_n306), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n314), .B1(new_n707), .B2(new_n694), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n624), .B2(new_n626), .ZN(new_n709));
  INV_X1    g523(.A(new_n504), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n573), .A3(new_n710), .A4(new_n647), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  AOI21_X1  g526(.A(new_n502), .B1(new_n624), .B2(new_n626), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n528), .A2(new_n529), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n533), .B1(new_n522), .B2(new_n527), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n526), .B1(new_n545), .B2(new_n537), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n507), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n609), .B2(G472), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n719), .A2(new_n605), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n713), .A2(new_n720), .A3(new_n669), .A4(new_n696), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR2_X1   g536(.A1(new_n623), .A2(new_n652), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n646), .B(new_n718), .C1(new_n609), .C2(G472), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n659), .A2(new_n723), .A3(new_n724), .A4(new_n696), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NAND2_X1  g540(.A1(new_n568), .A2(new_n508), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n553), .A3(new_n564), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n393), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n389), .B2(new_n392), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n289), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n284), .A2(new_n734), .A3(new_n288), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(G469), .A3(new_n293), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n300), .A2(new_n295), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n307), .B2(new_n300), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n313), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n732), .A2(new_n739), .A3(new_n605), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n723), .A4(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n740), .B(new_n723), .C1(new_n655), .C2(new_n656), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT110), .B(new_n741), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT111), .B(G131), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G33));
  NAND3_X1  g567(.A1(new_n573), .A2(new_n654), .A3(new_n740), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(new_n732), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n453), .A2(new_n622), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT43), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n453), .A2(new_n759), .A3(new_n622), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n647), .C1(new_n613), .C2(new_n614), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n300), .B1(new_n294), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n733), .A2(KEYINPUT45), .A3(new_n293), .A4(new_n735), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n737), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n308), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n314), .B(new_n671), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n764), .B(new_n772), .C1(new_n763), .C2(new_n762), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  OAI21_X1  g588(.A(new_n314), .B1(new_n769), .B2(new_n770), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n723), .A2(new_n628), .A3(new_n732), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n573), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NAND3_X1  g597(.A1(new_n605), .A2(new_n314), .A3(new_n393), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n668), .A2(new_n757), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n681), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n693), .A2(new_n695), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT49), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n758), .A2(new_n499), .A3(new_n760), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n731), .A3(new_n667), .A4(new_n666), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n720), .A2(new_n696), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT50), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n696), .A2(new_n732), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n786), .A2(new_n605), .A3(new_n797), .A4(new_n499), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n798), .A2(new_n452), .A3(new_n622), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n791), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n724), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n795), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n787), .A2(new_n313), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n777), .A2(new_n778), .A3(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n791), .A2(new_n720), .A3(new_n732), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n790), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n730), .A2(new_n605), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n810), .A2(new_n800), .A3(KEYINPUT115), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT115), .B1(new_n810), .B2(new_n800), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT48), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n798), .A2(new_n623), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n709), .A2(new_n791), .A3(new_n720), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n815), .A2(new_n495), .A3(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n809), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n803), .A2(new_n790), .A3(new_n808), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n725), .B1(new_n657), .B2(new_n660), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n689), .B2(new_n686), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n659), .A2(new_n669), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n647), .A2(new_n652), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n681), .A3(new_n739), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n659), .A2(new_n723), .A3(new_n696), .A4(new_n724), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n646), .B(new_n653), .C1(new_n567), .C2(new_n572), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(new_n687), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n690), .A2(new_n829), .A3(KEYINPUT52), .A4(new_n825), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n697), .A2(new_n701), .A3(new_n711), .A4(new_n721), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n452), .A2(new_n493), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n452), .B2(new_n622), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n394), .A3(new_n502), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n615), .A2(new_n836), .A3(new_n629), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n648), .A2(new_n837), .A3(new_n606), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n636), .A2(new_n637), .ZN(new_n839));
  INV_X1    g653(.A(new_n652), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n451), .A2(new_n493), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n839), .A2(new_n841), .A3(new_n646), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n573), .A2(new_n658), .A3(new_n732), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n724), .A2(new_n723), .A3(new_n732), .A4(new_n739), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n754), .A3(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n833), .A2(new_n838), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n749), .A3(new_n750), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT53), .B1(new_n832), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n846), .A2(new_n749), .A3(KEYINPUT112), .A4(new_n750), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n690), .A2(new_n829), .A3(new_n825), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(KEYINPUT113), .A3(new_n830), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n830), .A2(KEYINPUT113), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT54), .B(new_n848), .C1(new_n852), .C2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n857), .B1(new_n832), .B2(new_n847), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT114), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n833), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n845), .A2(new_n857), .ZN(new_n864));
  INV_X1    g678(.A(new_n838), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n747), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n856), .A2(new_n858), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n814), .A2(new_n817), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT116), .A2(new_n871), .A3(new_n819), .A4(new_n809), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n820), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n789), .B1(new_n873), .B2(new_n874), .ZN(G75));
  OR2_X1    g689(.A1(new_n384), .A2(new_n385), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT117), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT55), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n378), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n295), .B(new_n318), .C1(new_n861), .C2(new_n867), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(KEYINPUT56), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n286), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n880), .A2(KEYINPUT56), .A3(new_n879), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(G51));
  NAND2_X1  g700(.A1(new_n305), .A2(new_n306), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n861), .A2(new_n867), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n869), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n737), .B(KEYINPUT57), .Z(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n766), .A2(new_n767), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT118), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n888), .A2(G902), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n882), .B1(new_n893), .B2(new_n896), .ZN(G54));
  AND4_X1   g711(.A1(KEYINPUT58), .A2(new_n888), .A3(G475), .A4(G902), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n883), .B1(new_n898), .B2(new_n440), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n440), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n440), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G60));
  NOR2_X1   g718(.A1(new_n454), .A2(new_n295), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n621), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n882), .B1(new_n890), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n621), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n860), .B2(new_n869), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n908), .B(KEYINPUT120), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n912));
  INV_X1    g726(.A(new_n906), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n870), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n861), .A2(new_n868), .A3(new_n867), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n868), .B1(new_n861), .B2(new_n867), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n883), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n911), .A2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n888), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(new_n644), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n601), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n883), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n883), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  NOR2_X1   g744(.A1(new_n833), .A2(new_n838), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT121), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n286), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT122), .Z(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n501), .B2(new_n328), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(G898), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n877), .B1(new_n937), .B2(G953), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n938), .A3(new_n935), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G69));
  OAI21_X1  g756(.A(new_n517), .B1(new_n521), .B2(KEYINPUT30), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT123), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n434), .ZN(new_n945));
  NAND2_X1  g759(.A1(G900), .A2(G953), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n772), .A2(new_n605), .A3(new_n730), .A4(new_n823), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n773), .A2(new_n754), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n782), .A2(new_n822), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n751), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n945), .B(new_n946), .C1(new_n950), .C2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n822), .A2(new_n682), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n672), .A2(new_n756), .A3(new_n835), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n573), .A3(new_n605), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n773), .A2(new_n782), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n957), .A4(new_n954), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n951), .B1(new_n962), .B2(new_n945), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n286), .B1(G227), .B2(G900), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n951), .B2(KEYINPUT125), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n963), .B(new_n965), .Z(G72));
  XNOR2_X1  g780(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n960), .A2(new_n961), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n932), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n675), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n561), .A2(KEYINPUT127), .ZN(new_n974));
  AOI22_X1  g788(.A1(new_n561), .A2(KEYINPUT127), .B1(new_n522), .B2(new_n527), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n848), .B(new_n976), .C1(new_n852), .C2(new_n859), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n970), .B1(new_n950), .B2(new_n932), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n560), .A2(new_n536), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n882), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n973), .A2(new_n977), .A3(new_n980), .ZN(G57));
endmodule


