//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  AOI21_X1  g003(.A(KEYINPUT72), .B1(new_n189), .B2(G119), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n192), .B1(new_n191), .B2(new_n190), .ZN(new_n193));
  INV_X1    g007(.A(G110), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n188), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n199), .A2(KEYINPUT73), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(KEYINPUT73), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n209));
  XOR2_X1   g023(.A(new_n209), .B(KEYINPUT74), .Z(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(new_n206), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n208), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  OAI221_X1 g030(.A(new_n216), .B1(new_n193), .B2(new_n194), .C1(new_n197), .C2(new_n198), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  INV_X1    g033(.A(G221), .ZN(new_n220));
  INV_X1    g034(.A(G234), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n220), .A2(new_n221), .A3(G953), .ZN(new_n222));
  XOR2_X1   g036(.A(new_n219), .B(new_n222), .Z(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(new_n217), .A3(new_n223), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G217), .B1(new_n221), .B2(G902), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT71), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G902), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n225), .A2(new_n234), .A3(new_n226), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n225), .A2(new_n226), .A3(new_n237), .A4(new_n234), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n238), .A3(new_n229), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n227), .A2(KEYINPUT75), .A3(new_n230), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n233), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n242));
  NOR2_X1   g056(.A1(G237), .A2(G953), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G210), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n242), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G137), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n249), .A2(G137), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n249), .B2(G137), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT11), .A3(G134), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n250), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n211), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n262), .C2(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT64), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n261), .A3(new_n263), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n260), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n255), .A2(new_n257), .A3(new_n250), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n259), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n264), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(G143), .B(G146), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n272), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n284));
  INV_X1    g098(.A(G113), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT65), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(KEYINPUT2), .B2(G113), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n286), .A2(new_n288), .B1(KEYINPUT2), .B2(G113), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(G119), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n187), .B2(G116), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(KEYINPUT66), .A3(G119), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n289), .A2(new_n295), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT67), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n286), .A2(new_n288), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT2), .A2(G113), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n289), .A2(new_n295), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n283), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n259), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT68), .B1(new_n274), .B2(new_n259), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n271), .B1(new_n312), .B2(new_n281), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT67), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n309), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n275), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n259), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n281), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n272), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT28), .A3(new_n307), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n248), .B(new_n308), .C1(new_n317), .C2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(KEYINPUT30), .A3(new_n272), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  INV_X1    g140(.A(new_n282), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n271), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n328), .A3(new_n307), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n316), .A2(new_n321), .A3(new_n272), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n247), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n313), .A2(new_n316), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(KEYINPUT28), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n313), .A2(new_n309), .A3(new_n316), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n247), .A2(new_n333), .ZN(new_n339));
  AOI21_X1  g153(.A(G902), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G472), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(KEYINPUT70), .A3(G472), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(new_n248), .A3(new_n330), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT31), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT31), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n329), .A2(new_n349), .A3(new_n248), .A4(new_n330), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n336), .A2(new_n337), .B1(new_n307), .B2(new_n283), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n348), .B(new_n350), .C1(new_n351), .C2(new_n248), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT32), .B1(new_n352), .B2(new_n353), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n241), .B1(new_n346), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT9), .B(G234), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n220), .B1(new_n360), .B2(new_n234), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n362), .B2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G101), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n363), .A2(new_n366), .A3(new_n370), .A4(new_n367), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(KEYINPUT4), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n373), .A3(G101), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n281), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n365), .A2(G104), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n379));
  XNOR2_X1  g193(.A(G104), .B(G107), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n378), .A2(new_n381), .B1(new_n382), .B2(new_n370), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n268), .A2(new_n270), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT10), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n189), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n270), .B1(new_n386), .B2(new_n278), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n388));
  AOI211_X1 g202(.A(new_n379), .B(new_n370), .C1(new_n376), .C2(new_n367), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n387), .B(new_n371), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n375), .B(new_n385), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT78), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n385), .A2(new_n375), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n397), .B(new_n398), .C1(new_n394), .C2(new_n393), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n312), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G140), .ZN(new_n401));
  INV_X1    g215(.A(G227), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n401), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n385), .A2(new_n375), .ZN(new_n405));
  INV_X1    g219(.A(new_n394), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n319), .A2(new_n320), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT12), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n390), .B1(new_n383), .B2(new_n384), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n395), .A2(new_n312), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n404), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n420), .A2(KEYINPUT79), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n423));
  INV_X1    g237(.A(new_n404), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n395), .B2(new_n312), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n409), .B1(new_n395), .B2(KEYINPUT78), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n399), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n408), .A2(new_n409), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n415), .A2(new_n416), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n234), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n423), .B1(new_n431), .B2(G469), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n422), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n410), .A2(new_n429), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n424), .B1(new_n400), .B2(new_n428), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n418), .B1(new_n426), .B2(new_n399), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n438), .A2(KEYINPUT80), .A3(new_n424), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n421), .B(new_n234), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n361), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT81), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n285), .B1(new_n291), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n299), .B2(new_n446), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n383), .A2(new_n448), .A3(new_n305), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n372), .A2(new_n374), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n445), .B(new_n449), .C1(new_n316), .C2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n298), .B2(new_n306), .ZN(new_n452));
  INV_X1    g266(.A(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n444), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n454), .A3(KEYINPUT6), .ZN(new_n455));
  AOI21_X1  g269(.A(G125), .B1(new_n268), .B2(new_n270), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n205), .B1(new_n277), .B2(new_n280), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G953), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G224), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n460), .B(KEYINPUT82), .Z(new_n461));
  XNOR2_X1  g275(.A(new_n458), .B(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n444), .C1(new_n452), .C2(new_n453), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(KEYINPUT84), .A3(G224), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n460), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n466), .B(new_n469), .C1(new_n456), .C2(new_n457), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n460), .B1(new_n471), .B2(KEYINPUT7), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n471), .B2(KEYINPUT7), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n458), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n444), .B(KEYINPUT8), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n448), .A2(new_n305), .ZN(new_n476));
  INV_X1    g290(.A(new_n383), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n449), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n480), .B2(new_n451), .ZN(new_n481));
  OAI21_X1  g295(.A(G210), .B1(G237), .B2(G902), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n465), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n482), .B(KEYINPUT85), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n465), .B2(new_n481), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n442), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n442), .C1(new_n483), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n492));
  INV_X1    g306(.A(new_n209), .ZN(new_n493));
  AOI21_X1  g307(.A(G146), .B1(new_n207), .B2(new_n208), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n215), .A2(KEYINPUT93), .A3(new_n209), .ZN(new_n496));
  INV_X1    g310(.A(G237), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n459), .A3(G214), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n243), .B(G214), .C1(new_n499), .C2(G143), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT17), .A3(G131), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT94), .A4(new_n504), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n503), .B2(G131), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT92), .A4(new_n258), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n503), .A2(G131), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n507), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n362), .ZN(new_n518));
  NAND2_X1  g332(.A1(KEYINPUT18), .A2(G131), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n501), .B2(new_n502), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n522), .B(new_n519), .C1(new_n501), .C2(new_n502), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n204), .A2(new_n206), .A3(new_n211), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n211), .B1(new_n204), .B2(new_n206), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n204), .A2(new_n206), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G146), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT90), .A3(new_n212), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n501), .A2(new_n502), .A3(new_n519), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT91), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n520), .B(KEYINPUT89), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n516), .A2(new_n518), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n518), .B1(new_n516), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n234), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G475), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n529), .B(KEYINPUT19), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n210), .B(new_n546), .C1(G146), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n518), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n516), .A2(new_n518), .A3(new_n539), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n545), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI211_X1 g369(.A(KEYINPUT20), .B(new_n545), .C1(new_n551), .C2(new_n552), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n543), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n360), .A2(G217), .A3(new_n459), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n262), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n189), .A2(G143), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n249), .ZN(new_n562));
  XNOR2_X1  g376(.A(G116), .B(G122), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n365), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n365), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n560), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT13), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n262), .A2(G128), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n560), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT95), .B1(new_n560), .B2(new_n572), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n567), .B1(G134), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n562), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n249), .B1(new_n560), .B2(new_n561), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n564), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n290), .A2(KEYINPUT14), .A3(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G107), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT14), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n563), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n559), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n559), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n575), .A2(G134), .ZN(new_n587));
  OAI221_X1 g401(.A(new_n586), .B1(new_n583), .B2(new_n579), .C1(new_n587), .C2(new_n567), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n558), .B1(new_n589), .B2(new_n234), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT96), .B(G902), .C1(new_n585), .C2(new_n588), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n459), .A2(G952), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(G234), .B2(G237), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n234), .B(new_n459), .C1(G234), .C2(G237), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT21), .B(G898), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n557), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n358), .A2(new_n441), .A3(new_n491), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n431), .A2(G469), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n431), .A2(new_n423), .A3(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n440), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n241), .ZN(new_n610));
  INV_X1    g424(.A(new_n361), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n352), .A2(new_n234), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n612), .A2(G472), .B1(new_n353), .B2(new_n352), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n234), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n591), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(new_n618), .A3(new_n591), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n589), .B(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(G478), .A3(new_n234), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n557), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n482), .B1(new_n465), .B2(new_n481), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n483), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n602), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n442), .A3(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n614), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT34), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  INV_X1    g445(.A(new_n554), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n518), .B1(new_n539), .B2(new_n548), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n505), .A2(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n634), .A2(new_n508), .B1(new_n538), .B2(new_n534), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n518), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n632), .B1(new_n636), .B2(new_n545), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n553), .A2(new_n554), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(KEYINPUT98), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n595), .A2(new_n593), .B1(new_n542), .B2(G475), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n553), .A2(new_n641), .A3(new_n554), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n614), .A2(new_n628), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NAND3_X1  g460(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n213), .B2(new_n217), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n213), .A2(new_n648), .A3(new_n217), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n650), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n230), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n239), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n491), .A2(new_n603), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  OAI211_X1 g474(.A(new_n656), .B(new_n442), .C1(new_n483), .C2(new_n625), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n346), .B2(new_n357), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n600), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n599), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n639), .A2(new_n640), .A3(new_n642), .A4(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT100), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT100), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n662), .A2(new_n441), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XNOR2_X1  g485(.A(new_n666), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n441), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n330), .A2(new_n247), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n234), .B1(new_n676), .B2(new_n335), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n247), .B1(new_n329), .B2(new_n330), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n357), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT101), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n465), .A2(new_n481), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n484), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n465), .A2(new_n481), .A3(new_n482), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT38), .ZN(new_n686));
  INV_X1    g500(.A(new_n656), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT20), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n553), .A2(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n637), .A2(new_n689), .B1(G475), .B2(new_n542), .ZN(new_n690));
  INV_X1    g504(.A(new_n442), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n690), .A2(new_n691), .A3(new_n596), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n686), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n674), .A2(new_n675), .A3(new_n681), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND3_X1  g509(.A1(new_n557), .A2(new_n623), .A3(new_n666), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n662), .A2(new_n441), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(new_n440), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n400), .A2(new_n428), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n436), .A3(new_n404), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT80), .B1(new_n438), .B2(new_n424), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n434), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n421), .B1(new_n704), .B2(new_n234), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n700), .A2(new_n705), .A3(new_n361), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n628), .A2(new_n624), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n358), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT102), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n706), .A2(new_n358), .A3(new_n710), .A4(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NOR2_X1   g528(.A1(new_n628), .A2(new_n643), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n358), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND3_X1  g531(.A1(new_n706), .A2(new_n662), .A3(new_n603), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NOR2_X1   g533(.A1(new_n596), .A2(new_n691), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n626), .A3(new_n557), .A4(new_n627), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n612), .A2(G472), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n348), .A2(new_n350), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n338), .A2(new_n248), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n353), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n610), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n706), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NOR2_X1   g543(.A1(new_n700), .A2(new_n705), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n656), .A3(new_n725), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n696), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n626), .A2(new_n442), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n732), .A3(new_n611), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n440), .A2(new_n606), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n683), .A2(new_n442), .A3(new_n684), .A4(new_n611), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI211_X1 g554(.A(KEYINPUT103), .B(new_n738), .C1(new_n440), .C2(new_n606), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n358), .B(new_n697), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n739), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n737), .A2(new_n736), .A3(new_n739), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n557), .A2(KEYINPUT42), .A3(new_n623), .A4(new_n666), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n355), .B1(new_n344), .B2(new_n345), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n356), .A2(KEYINPUT105), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n751), .B(KEYINPUT32), .C1(new_n352), .C2(new_n353), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n241), .B(new_n748), .C1(new_n749), .C2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n742), .A2(new_n743), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n258), .ZN(G33));
  INV_X1    g570(.A(KEYINPUT100), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n667), .B(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(new_n358), .C1(new_n740), .C2(new_n741), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT106), .B(G134), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G36));
  AND2_X1   g575(.A1(new_n620), .A2(new_n622), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n557), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n613), .A3(new_n687), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n683), .A2(new_n442), .A3(new_n684), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n427), .A2(new_n430), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n772), .B2(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(KEYINPUT45), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n421), .A2(new_n234), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n440), .B1(new_n776), .B2(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT107), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n361), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n672), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT108), .A3(new_n672), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n771), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n256), .ZN(G39));
  NAND2_X1  g602(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(new_n789), .ZN(new_n792));
  OAI22_X1  g606(.A1(new_n781), .A2(new_n361), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n346), .A2(new_n357), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n794), .A2(new_n610), .A3(new_n696), .A4(new_n768), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT110), .B(G140), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G42));
  NAND4_X1  g612(.A1(new_n763), .A2(new_n610), .A3(new_n442), .A4(new_n611), .ZN(new_n799));
  INV_X1    g613(.A(new_n730), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(KEYINPUT49), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT111), .Z(new_n802));
  INV_X1    g616(.A(new_n686), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n800), .B2(KEYINPUT49), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n802), .A2(new_n681), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n706), .A2(new_n769), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n765), .A2(new_n665), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n749), .A2(new_n753), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n610), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n681), .A2(new_n241), .A3(new_n665), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n807), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n624), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n765), .A2(new_n665), .A3(new_n726), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n706), .A2(new_n733), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n813), .A2(new_n598), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n706), .A2(new_n691), .A3(new_n803), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(KEYINPUT50), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT50), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n790), .A2(new_n793), .B1(new_n361), .B2(new_n730), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n817), .A2(new_n768), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n690), .A2(new_n762), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n815), .A2(new_n831), .B1(new_n731), .B2(new_n809), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT118), .Z(new_n833));
  OAI21_X1  g647(.A(new_n820), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n732), .B1(new_n740), .B2(new_n741), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n656), .A2(new_n543), .A3(new_n596), .A4(new_n666), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n639), .A2(new_n642), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n836), .A2(new_n837), .A3(new_n768), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n441), .A2(new_n794), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n759), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n755), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n690), .B2(new_n762), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n557), .A2(KEYINPUT112), .A3(new_n623), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n690), .A2(new_n597), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n602), .B1(new_n488), .B2(new_n490), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(new_n614), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT113), .A3(new_n604), .A4(new_n658), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n609), .A2(new_n491), .A3(new_n603), .A4(new_n611), .ZN(new_n852));
  INV_X1    g666(.A(new_n345), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT70), .B1(new_n341), .B2(G472), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n356), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n354), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n610), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n852), .A2(new_n858), .B1(new_n647), .B2(new_n657), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n848), .A2(new_n614), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n850), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n716), .A2(new_n718), .A3(new_n728), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n711), .B2(new_n709), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n841), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n239), .A2(new_n655), .A3(new_n611), .A4(new_n666), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n557), .A2(new_n867), .A3(new_n626), .A4(new_n720), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n680), .A3(new_n737), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n670), .A2(new_n698), .A3(new_n734), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n441), .B(new_n662), .C1(new_n758), .C2(new_n697), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT52), .A3(new_n734), .A4(new_n869), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT53), .A4(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n870), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(new_n870), .B2(KEYINPUT114), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n865), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n875), .A2(new_n841), .A3(new_n862), .A4(new_n864), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT115), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT54), .B(new_n876), .C1(new_n880), .C2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n716), .A2(new_n718), .A3(new_n728), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n712), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n861), .B2(new_n850), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n879), .A3(KEYINPUT53), .A4(new_n841), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n881), .A2(new_n882), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT116), .A4(new_n890), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n884), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n827), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(KEYINPUT117), .A3(new_n828), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n832), .B1(new_n824), .B2(new_n825), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n827), .B2(new_n829), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n834), .B(new_n895), .C1(new_n821), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n805), .B1(new_n902), .B2(new_n903), .ZN(G75));
  NOR2_X1   g718(.A1(new_n459), .A2(G952), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT119), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n455), .A2(new_n464), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n462), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n234), .B1(new_n888), .B2(new_n889), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G210), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n484), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n910), .A2(new_n913), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n907), .B(new_n914), .C1(new_n915), .C2(new_n916), .ZN(G51));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n774), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n704), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n888), .A2(new_n889), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n891), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n775), .B(KEYINPUT57), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n920), .B1(KEYINPUT120), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n926), .A2(KEYINPUT120), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n905), .B1(new_n927), .B2(new_n928), .ZN(G54));
  AND3_X1   g743(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  INV_X1    g744(.A(new_n636), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n905), .ZN(G60));
  XNOR2_X1  g748(.A(new_n621), .B(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT123), .B1(new_n924), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n890), .B1(new_n888), .B2(new_n889), .ZN(new_n942));
  OAI211_X1 g756(.A(KEYINPUT123), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n906), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n895), .B2(new_n938), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT124), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n946), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n907), .B1(new_n951), .B2(new_n943), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n948), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n947), .A2(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n888), .B2(new_n889), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n653), .B2(new_n654), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n959), .B(new_n906), .C1(new_n227), .C2(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G66));
  INV_X1    g777(.A(new_n601), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n459), .B1(new_n964), .B2(G224), .ZN(new_n965));
  INV_X1    g779(.A(new_n887), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n459), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n908), .B1(G898), .B2(new_n459), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(G69));
  AND2_X1   g783(.A1(new_n873), .A2(new_n734), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT62), .B1(new_n694), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n694), .A2(KEYINPUT62), .A3(new_n970), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n796), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n358), .A2(new_n769), .A3(new_n846), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n673), .ZN(new_n975));
  NOR4_X1   g789(.A1(new_n973), .A2(new_n787), .A3(G953), .A4(new_n975), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n402), .A2(new_n663), .A3(new_n459), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n325), .A2(new_n328), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n547), .ZN(new_n979));
  OR3_X1    g793(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n771), .ZN(new_n981));
  INV_X1    g795(.A(new_n786), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT108), .B1(new_n782), .B2(new_n672), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n984), .A2(KEYINPUT126), .A3(new_n970), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT126), .B1(new_n984), .B2(new_n970), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n692), .A2(new_n626), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n988), .B(new_n811), .C1(new_n785), .C2(new_n786), .ZN(new_n989));
  INV_X1    g803(.A(new_n755), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n796), .A2(new_n990), .A3(new_n759), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(G953), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n402), .A2(G900), .A3(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n979), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n980), .B1(new_n993), .B2(new_n995), .ZN(G72));
  OAI211_X1 g810(.A(new_n992), .B(new_n887), .C1(new_n985), .C2(new_n986), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT63), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n331), .A2(new_n248), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1002), .A2(new_n678), .A3(new_n999), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n876), .B(new_n1004), .C1(new_n880), .C2(new_n883), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n984), .B(new_n887), .C1(new_n673), .C2(new_n974), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1000), .B1(new_n1006), .B2(new_n973), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n905), .B1(new_n1007), .B2(new_n678), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1003), .A2(new_n1005), .A3(new_n1008), .ZN(G57));
endmodule


