

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721;

  XNOR2_X1 U364 ( .A(n689), .B(n688), .ZN(n343) );
  XNOR2_X2 U365 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X2 U366 ( .A(n360), .B(n412), .ZN(n359) );
  XNOR2_X2 U367 ( .A(n488), .B(KEYINPUT16), .ZN(n366) );
  NOR2_X1 U368 ( .A1(n343), .A2(n691), .ZN(G66) );
  XNOR2_X2 U369 ( .A(n692), .B(KEYINPUT70), .ZN(n367) );
  INV_X1 U370 ( .A(G953), .ZN(n710) );
  BUF_X1 U371 ( .A(G107), .Z(n344) );
  AND2_X2 U372 ( .A1(n362), .A2(n361), .ZN(n351) );
  NAND2_X2 U373 ( .A1(n401), .A2(n403), .ZN(n400) );
  AND2_X2 U374 ( .A1(n591), .A2(n450), .ZN(n401) );
  NOR2_X2 U375 ( .A1(n709), .A2(KEYINPUT2), .ZN(n403) );
  XNOR2_X2 U376 ( .A(n367), .B(n466), .ZN(n432) );
  XNOR2_X2 U377 ( .A(n565), .B(KEYINPUT1), .ZN(n508) );
  INV_X1 U378 ( .A(n696), .ZN(n591) );
  XNOR2_X1 U379 ( .A(n419), .B(n418), .ZN(n542) );
  NAND2_X1 U380 ( .A1(n402), .A2(n399), .ZN(n398) );
  XNOR2_X1 U381 ( .A(n590), .B(KEYINPUT78), .ZN(n709) );
  AND2_X1 U382 ( .A1(n511), .A2(n721), .ZN(n347) );
  NAND2_X1 U383 ( .A1(n508), .A2(n458), .ZN(n519) );
  XNOR2_X1 U384 ( .A(n443), .B(n444), .ZN(n705) );
  XNOR2_X1 U385 ( .A(KEYINPUT94), .B(G146), .ZN(n429) );
  XNOR2_X1 U386 ( .A(G143), .B(G128), .ZN(n433) );
  XNOR2_X1 U387 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n706) );
  XNOR2_X2 U388 ( .A(n345), .B(n437), .ZN(n565) );
  NAND2_X1 U389 ( .A1(n683), .A2(n496), .ZN(n345) );
  XNOR2_X1 U390 ( .A(n542), .B(KEYINPUT19), .ZN(n570) );
  XNOR2_X1 U391 ( .A(n569), .B(KEYINPUT46), .ZN(n350) );
  BUF_X1 U392 ( .A(n363), .Z(n346) );
  XNOR2_X1 U393 ( .A(n505), .B(KEYINPUT22), .ZN(n363) );
  NAND2_X1 U394 ( .A1(n511), .A2(n721), .ZN(n530) );
  NOR2_X1 U395 ( .A1(n521), .A2(n504), .ZN(n505) );
  XNOR2_X2 U396 ( .A(n369), .B(n499), .ZN(n506) );
  XNOR2_X2 U397 ( .A(n385), .B(n354), .ZN(n696) );
  XNOR2_X2 U398 ( .A(G146), .B(G125), .ZN(n443) );
  INV_X1 U399 ( .A(KEYINPUT84), .ZN(n418) );
  XNOR2_X1 U400 ( .A(n353), .B(n453), .ZN(n538) );
  XNOR2_X1 U401 ( .A(n594), .B(n355), .ZN(n599) );
  XNOR2_X1 U402 ( .A(n404), .B(n410), .ZN(n411) );
  INV_X1 U403 ( .A(KEYINPUT48), .ZN(n379) );
  NAND2_X1 U404 ( .A1(n381), .A2(KEYINPUT48), .ZN(n380) );
  NAND2_X1 U405 ( .A1(G234), .A2(G237), .ZN(n420) );
  INV_X1 U406 ( .A(KEYINPUT44), .ZN(n387) );
  XNOR2_X1 U407 ( .A(n397), .B(G119), .ZN(n396) );
  INV_X1 U408 ( .A(KEYINPUT3), .ZN(n397) );
  XNOR2_X1 U409 ( .A(G143), .B(G131), .ZN(n478) );
  INV_X1 U410 ( .A(G140), .ZN(n477) );
  XNOR2_X1 U411 ( .A(G113), .B(G104), .ZN(n481) );
  XOR2_X1 U412 ( .A(KEYINPUT12), .B(G122), .Z(n482) );
  XOR2_X1 U413 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n475) );
  NOR2_X1 U414 ( .A1(n592), .A2(n547), .ZN(n548) );
  XNOR2_X1 U415 ( .A(n440), .B(KEYINPUT23), .ZN(n441) );
  INV_X1 U416 ( .A(G119), .ZN(n440) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(G140), .ZN(n442) );
  XNOR2_X1 U418 ( .A(G137), .B(G128), .ZN(n438) );
  XOR2_X1 U419 ( .A(KEYINPUT24), .B(G110), .Z(n439) );
  XNOR2_X1 U420 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n444) );
  XNOR2_X1 U421 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n446) );
  XNOR2_X1 U422 ( .A(n556), .B(n555), .ZN(n586) );
  NOR2_X1 U423 ( .A1(n570), .A2(n425), .ZN(n427) );
  NAND2_X1 U424 ( .A1(n393), .A2(n391), .ZN(n373) );
  AND2_X1 U425 ( .A1(n405), .A2(n596), .ZN(n368) );
  XNOR2_X1 U426 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n355) );
  XOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT90), .Z(n409) );
  XOR2_X1 U428 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n408) );
  XNOR2_X1 U429 ( .A(n605), .B(KEYINPUT51), .ZN(n356) );
  NOR2_X1 U430 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U431 ( .A1(G953), .A2(G237), .ZN(n474) );
  XNOR2_X1 U432 ( .A(n411), .B(n414), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n358), .B(n432), .ZN(n364) );
  INV_X1 U434 ( .A(n443), .ZN(n414) );
  XOR2_X1 U435 ( .A(KEYINPUT38), .B(n573), .Z(n607) );
  BUF_X1 U436 ( .A(n553), .Z(n573) );
  XNOR2_X1 U437 ( .A(G137), .B(G131), .ZN(n434) );
  NAND2_X1 U438 ( .A1(n347), .A2(n387), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U440 ( .A1(n624), .A2(n623), .ZN(n625) );
  AND2_X1 U441 ( .A1(n548), .A2(n565), .ZN(n549) );
  NAND2_X1 U442 ( .A1(n538), .A2(n502), .ZN(n592) );
  XNOR2_X1 U443 ( .A(n448), .B(n382), .ZN(n688) );
  XNOR2_X1 U444 ( .A(n352), .B(n449), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n442), .B(n441), .ZN(n445) );
  XNOR2_X1 U446 ( .A(n633), .B(KEYINPUT88), .ZN(n676) );
  XNOR2_X1 U447 ( .A(n559), .B(n558), .ZN(n719) );
  XNOR2_X1 U448 ( .A(KEYINPUT112), .B(KEYINPUT36), .ZN(n544) );
  AND2_X1 U449 ( .A1(n510), .A2(n596), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n357), .B(KEYINPUT121), .ZN(n371) );
  INV_X1 U451 ( .A(n507), .ZN(n654) );
  NAND2_X1 U452 ( .A1(n578), .A2(n577), .ZN(n348) );
  NOR2_X1 U453 ( .A1(n523), .A2(n525), .ZN(n349) );
  AND2_X1 U454 ( .A1(G221), .A2(n491), .ZN(n352) );
  NOR2_X1 U455 ( .A1(n688), .A2(G902), .ZN(n353) );
  INV_X1 U456 ( .A(n348), .ZN(n381) );
  XNOR2_X1 U457 ( .A(KEYINPUT79), .B(KEYINPUT45), .ZN(n354) );
  XNOR2_X1 U458 ( .A(n364), .B(n365), .ZN(n671) );
  NOR2_X1 U459 ( .A1(n356), .A2(n622), .ZN(n617) );
  NAND2_X1 U460 ( .A1(n373), .A2(n372), .ZN(n357) );
  NAND2_X1 U461 ( .A1(n394), .A2(n591), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n358), .B(n693), .ZN(n695) );
  XNOR2_X2 U463 ( .A(n366), .B(n462), .ZN(n358) );
  XNOR2_X2 U464 ( .A(n359), .B(n396), .ZN(n462) );
  XNOR2_X2 U465 ( .A(G113), .B(KEYINPUT89), .ZN(n360) );
  INV_X1 U466 ( .A(n528), .ZN(n361) );
  XNOR2_X1 U467 ( .A(n362), .B(G101), .ZN(n647) );
  NAND2_X1 U468 ( .A1(n515), .A2(n538), .ZN(n362) );
  NAND2_X1 U469 ( .A1(n363), .A2(n512), .ZN(n514) );
  NAND2_X1 U470 ( .A1(n363), .A2(n383), .ZN(n384) );
  NAND2_X1 U471 ( .A1(n346), .A2(n368), .ZN(n507) );
  AND2_X2 U472 ( .A1(n506), .A2(n507), .ZN(n511) );
  NAND2_X1 U473 ( .A1(n370), .A2(n349), .ZN(n369) );
  XNOR2_X1 U474 ( .A(n473), .B(KEYINPUT34), .ZN(n370) );
  NAND2_X1 U475 ( .A1(n371), .A2(n710), .ZN(n626) );
  NAND2_X1 U476 ( .A1(n403), .A2(n591), .ZN(n372) );
  NAND2_X1 U477 ( .A1(n374), .A2(n350), .ZN(n376) );
  NOR2_X1 U478 ( .A1(n666), .A2(n348), .ZN(n374) );
  NOR2_X2 U479 ( .A1(n546), .A2(n593), .ZN(n666) );
  NAND2_X1 U480 ( .A1(n375), .A2(n377), .ZN(n589) );
  NAND2_X1 U481 ( .A1(n376), .A2(n379), .ZN(n375) );
  NAND2_X1 U482 ( .A1(n378), .A2(n350), .ZN(n377) );
  NOR2_X1 U483 ( .A1(n666), .A2(n380), .ZN(n378) );
  XNOR2_X2 U484 ( .A(n384), .B(KEYINPUT32), .ZN(n721) );
  NAND2_X1 U485 ( .A1(n529), .A2(n351), .ZN(n389) );
  NAND2_X1 U486 ( .A1(n388), .A2(n386), .ZN(n385) );
  XNOR2_X1 U487 ( .A(n389), .B(KEYINPUT83), .ZN(n388) );
  XNOR2_X2 U488 ( .A(n390), .B(G110), .ZN(n692) );
  XNOR2_X2 U489 ( .A(G104), .B(KEYINPUT73), .ZN(n390) );
  OR2_X1 U490 ( .A1(n696), .A2(n590), .ZN(n402) );
  NAND2_X1 U491 ( .A1(n625), .A2(n392), .ZN(n391) );
  INV_X1 U492 ( .A(KEYINPUT2), .ZN(n392) );
  AND2_X1 U493 ( .A1(n625), .A2(n395), .ZN(n394) );
  INV_X1 U494 ( .A(n590), .ZN(n395) );
  NAND2_X2 U495 ( .A1(n400), .A2(n398), .ZN(n670) );
  NOR2_X1 U496 ( .A1(n627), .A2(n392), .ZN(n399) );
  XOR2_X1 U497 ( .A(n408), .B(n407), .Z(n404) );
  NOR2_X1 U498 ( .A1(n508), .A2(n601), .ZN(n405) );
  INV_X1 U499 ( .A(n717), .ZN(n577) );
  INV_X1 U500 ( .A(n661), .ZN(n539) );
  XNOR2_X1 U501 ( .A(G116), .B(KEYINPUT72), .ZN(n465) );
  XNOR2_X1 U502 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U503 ( .A(n480), .B(n479), .ZN(n485) );
  INV_X1 U504 ( .A(KEYINPUT104), .ZN(n531) );
  INV_X1 U505 ( .A(KEYINPUT40), .ZN(n558) );
  INV_X1 U506 ( .A(KEYINPUT15), .ZN(n406) );
  XNOR2_X1 U507 ( .A(n406), .B(G902), .ZN(n450) );
  XNOR2_X1 U508 ( .A(G101), .B(n706), .ZN(n466) );
  NAND2_X1 U509 ( .A1(G224), .A2(n710), .ZN(n407) );
  XOR2_X1 U510 ( .A(n409), .B(n433), .Z(n410) );
  INV_X1 U511 ( .A(KEYINPUT69), .ZN(n412) );
  XNOR2_X2 U512 ( .A(G116), .B(G107), .ZN(n413) );
  XNOR2_X2 U513 ( .A(n413), .B(G122), .ZN(n488) );
  NOR2_X2 U514 ( .A1(n450), .A2(n671), .ZN(n416) );
  OR2_X1 U515 ( .A1(G237), .A2(G902), .ZN(n417) );
  NAND2_X1 U516 ( .A1(G210), .A2(n417), .ZN(n415) );
  XNOR2_X2 U517 ( .A(n416), .B(n415), .ZN(n553) );
  NAND2_X1 U518 ( .A1(G214), .A2(n417), .ZN(n606) );
  NAND2_X1 U519 ( .A1(n553), .A2(n606), .ZN(n419) );
  XNOR2_X1 U520 ( .A(n420), .B(KEYINPUT14), .ZN(n422) );
  NAND2_X1 U521 ( .A1(n422), .A2(G952), .ZN(n619) );
  NOR2_X1 U522 ( .A1(G953), .A2(n619), .ZN(n535) );
  XNOR2_X1 U523 ( .A(G898), .B(KEYINPUT91), .ZN(n699) );
  NAND2_X1 U524 ( .A1(n699), .A2(G953), .ZN(n421) );
  XNOR2_X1 U525 ( .A(n421), .B(KEYINPUT92), .ZN(n694) );
  NAND2_X1 U526 ( .A1(G902), .A2(n422), .ZN(n532) );
  NOR2_X1 U527 ( .A1(n694), .A2(n532), .ZN(n423) );
  XOR2_X1 U528 ( .A(KEYINPUT93), .B(n423), .Z(n424) );
  NOR2_X1 U529 ( .A1(n535), .A2(n424), .ZN(n425) );
  INV_X1 U530 ( .A(KEYINPUT0), .ZN(n426) );
  XNOR2_X2 U531 ( .A(n427), .B(n426), .ZN(n521) );
  NAND2_X1 U532 ( .A1(n710), .A2(G227), .ZN(n428) );
  XNOR2_X1 U533 ( .A(n428), .B(n344), .ZN(n430) );
  XNOR2_X1 U534 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U535 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U536 ( .A(n433), .B(G134), .ZN(n492) );
  XNOR2_X1 U537 ( .A(n492), .B(n434), .ZN(n463) );
  INV_X1 U538 ( .A(n442), .ZN(n435) );
  XNOR2_X1 U539 ( .A(n463), .B(n435), .ZN(n708) );
  XNOR2_X1 U540 ( .A(n436), .B(n708), .ZN(n683) );
  INV_X1 U541 ( .A(G902), .ZN(n496) );
  XNOR2_X1 U542 ( .A(KEYINPUT68), .B(G469), .ZN(n437) );
  XNOR2_X1 U543 ( .A(n439), .B(n438), .ZN(n449) );
  XNOR2_X1 U544 ( .A(n445), .B(n705), .ZN(n448) );
  NAND2_X1 U545 ( .A1(n710), .A2(G234), .ZN(n447) );
  XNOR2_X1 U546 ( .A(n447), .B(n446), .ZN(n491) );
  INV_X1 U547 ( .A(n450), .ZN(n627) );
  NAND2_X1 U548 ( .A1(G234), .A2(n627), .ZN(n451) );
  XNOR2_X1 U549 ( .A(KEYINPUT20), .B(n451), .ZN(n454) );
  NAND2_X1 U550 ( .A1(G217), .A2(n454), .ZN(n452) );
  XNOR2_X1 U551 ( .A(n452), .B(KEYINPUT25), .ZN(n453) );
  XOR2_X1 U552 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n456) );
  NAND2_X1 U553 ( .A1(n454), .A2(G221), .ZN(n455) );
  XNOR2_X1 U554 ( .A(n456), .B(n455), .ZN(n595) );
  INV_X1 U555 ( .A(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n595), .B(n457), .ZN(n502) );
  INV_X1 U557 ( .A(n592), .ZN(n458) );
  XOR2_X1 U558 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n460) );
  NAND2_X1 U559 ( .A1(n474), .A2(G210), .ZN(n459) );
  XNOR2_X1 U560 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U561 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U562 ( .A(n464), .B(n463), .ZN(n469) );
  XOR2_X1 U563 ( .A(n467), .B(G146), .Z(n468) );
  XNOR2_X1 U564 ( .A(n469), .B(n468), .ZN(n629) );
  NAND2_X1 U565 ( .A1(n629), .A2(n496), .ZN(n471) );
  XOR2_X1 U566 ( .A(G472), .B(KEYINPUT71), .Z(n470) );
  XNOR2_X2 U567 ( .A(n471), .B(n470), .ZN(n601) );
  XNOR2_X1 U568 ( .A(n601), .B(KEYINPUT6), .ZN(n541) );
  NOR2_X1 U569 ( .A1(n519), .A2(n541), .ZN(n472) );
  XNOR2_X1 U570 ( .A(n472), .B(KEYINPUT33), .ZN(n621) );
  NOR2_X1 U571 ( .A1(n521), .A2(n621), .ZN(n473) );
  NAND2_X1 U572 ( .A1(G214), .A2(n474), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n476), .B(n475), .ZN(n480) );
  XOR2_X1 U574 ( .A(n482), .B(n481), .Z(n483) );
  XNOR2_X1 U575 ( .A(n483), .B(n705), .ZN(n484) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n637) );
  NAND2_X1 U577 ( .A1(n637), .A2(n496), .ZN(n487) );
  XNOR2_X1 U578 ( .A(KEYINPUT13), .B(G475), .ZN(n486) );
  XNOR2_X2 U579 ( .A(n487), .B(n486), .ZN(n523) );
  XOR2_X1 U580 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n490) );
  XNOR2_X1 U581 ( .A(n488), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U582 ( .A(n490), .B(n489), .ZN(n495) );
  NAND2_X1 U583 ( .A1(n491), .A2(G217), .ZN(n493) );
  XOR2_X1 U584 ( .A(n493), .B(n492), .Z(n494) );
  XNOR2_X1 U585 ( .A(n495), .B(n494), .ZN(n643) );
  NAND2_X1 U586 ( .A1(n643), .A2(n496), .ZN(n498) );
  INV_X1 U587 ( .A(G478), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n498), .B(n497), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT75), .B(KEYINPUT35), .ZN(n499) );
  XOR2_X1 U590 ( .A(G122), .B(KEYINPUT127), .Z(n500) );
  XNOR2_X1 U591 ( .A(n506), .B(n500), .ZN(G24) );
  NAND2_X1 U592 ( .A1(n525), .A2(n523), .ZN(n610) );
  INV_X1 U593 ( .A(n610), .ZN(n501) );
  NAND2_X1 U594 ( .A1(n502), .A2(n501), .ZN(n503) );
  XOR2_X1 U595 ( .A(KEYINPUT103), .B(n503), .Z(n504) );
  INV_X1 U596 ( .A(n538), .ZN(n596) );
  INV_X1 U597 ( .A(n508), .ZN(n593) );
  XOR2_X1 U598 ( .A(KEYINPUT76), .B(n541), .Z(n509) );
  NOR2_X1 U599 ( .A1(n593), .A2(n509), .ZN(n510) );
  NAND2_X1 U600 ( .A1(n530), .A2(KEYINPUT44), .ZN(n529) );
  AND2_X1 U601 ( .A1(n593), .A2(n541), .ZN(n512) );
  INV_X1 U602 ( .A(KEYINPUT82), .ZN(n513) );
  XNOR2_X1 U603 ( .A(n514), .B(n513), .ZN(n515) );
  NOR2_X1 U604 ( .A1(n601), .A2(n592), .ZN(n516) );
  NAND2_X1 U605 ( .A1(n516), .A2(n565), .ZN(n517) );
  OR2_X1 U606 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U607 ( .A(KEYINPUT98), .B(n518), .ZN(n650) );
  INV_X1 U608 ( .A(n519), .ZN(n520) );
  NAND2_X1 U609 ( .A1(n520), .A2(n601), .ZN(n603) );
  NOR2_X1 U610 ( .A1(n521), .A2(n603), .ZN(n522) );
  XNOR2_X1 U611 ( .A(n522), .B(KEYINPUT31), .ZN(n663) );
  AND2_X1 U612 ( .A1(n650), .A2(n663), .ZN(n527) );
  XOR2_X1 U613 ( .A(n523), .B(KEYINPUT100), .Z(n526) );
  AND2_X1 U614 ( .A1(n526), .A2(n525), .ZN(n524) );
  XNOR2_X1 U615 ( .A(KEYINPUT102), .B(n524), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n526), .A2(n525), .ZN(n649) );
  NOR2_X1 U617 ( .A1(n557), .A2(n649), .ZN(n612) );
  NOR2_X1 U618 ( .A1(n527), .A2(n612), .ZN(n528) );
  XNOR2_X1 U619 ( .A(n557), .B(n531), .ZN(n661) );
  OR2_X1 U620 ( .A1(n710), .A2(n532), .ZN(n533) );
  NOR2_X1 U621 ( .A1(G900), .A2(n533), .ZN(n534) );
  NOR2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n547) );
  NOR2_X1 U623 ( .A1(n547), .A2(n595), .ZN(n536) );
  XNOR2_X1 U624 ( .A(n536), .B(KEYINPUT67), .ZN(n537) );
  NOR2_X1 U625 ( .A1(n538), .A2(n537), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n539), .A2(n562), .ZN(n540) );
  NOR2_X1 U627 ( .A1(n541), .A2(n540), .ZN(n579) );
  XOR2_X1 U628 ( .A(n579), .B(KEYINPUT111), .Z(n543) );
  NAND2_X1 U629 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U630 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U631 ( .A(KEYINPUT81), .B(KEYINPUT39), .Z(n556) );
  XNOR2_X1 U632 ( .A(n549), .B(KEYINPUT74), .ZN(n552) );
  NAND2_X1 U633 ( .A1(n601), .A2(n606), .ZN(n550) );
  XOR2_X1 U634 ( .A(KEYINPUT30), .B(n550), .Z(n551) );
  NAND2_X1 U635 ( .A1(n552), .A2(n551), .ZN(n574) );
  INV_X1 U636 ( .A(n574), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n554), .A2(n607), .ZN(n555) );
  NAND2_X1 U638 ( .A1(n586), .A2(n557), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n607), .A2(n606), .ZN(n611) );
  NOR2_X1 U640 ( .A1(n611), .A2(n610), .ZN(n560) );
  XNOR2_X1 U641 ( .A(n560), .B(KEYINPUT41), .ZN(n622) );
  XOR2_X1 U642 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n561) );
  XNOR2_X1 U643 ( .A(KEYINPUT110), .B(n561), .ZN(n564) );
  NAND2_X1 U644 ( .A1(n562), .A2(n601), .ZN(n563) );
  XOR2_X1 U645 ( .A(n564), .B(n563), .Z(n567) );
  XNOR2_X1 U646 ( .A(n565), .B(KEYINPUT108), .ZN(n566) );
  NAND2_X1 U647 ( .A1(n567), .A2(n566), .ZN(n571) );
  NOR2_X1 U648 ( .A1(n622), .A2(n571), .ZN(n568) );
  XNOR2_X1 U649 ( .A(KEYINPUT42), .B(n568), .ZN(n718) );
  NOR2_X1 U650 ( .A1(n719), .A2(n718), .ZN(n569) );
  OR2_X1 U651 ( .A1(n571), .A2(n570), .ZN(n658) );
  NOR2_X1 U652 ( .A1(n658), .A2(n612), .ZN(n572) );
  XNOR2_X1 U653 ( .A(n572), .B(KEYINPUT47), .ZN(n578) );
  INV_X1 U654 ( .A(n573), .ZN(n583) );
  NOR2_X1 U655 ( .A1(n583), .A2(n574), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n349), .A2(n575), .ZN(n576) );
  XNOR2_X1 U657 ( .A(KEYINPUT107), .B(n576), .ZN(n717) );
  NAND2_X1 U658 ( .A1(n579), .A2(n606), .ZN(n580) );
  NOR2_X1 U659 ( .A1(n580), .A2(n508), .ZN(n582) );
  XNOR2_X1 U660 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n581) );
  XNOR2_X1 U661 ( .A(n582), .B(n581), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U663 ( .A(KEYINPUT106), .B(n585), .Z(n720) );
  NAND2_X1 U664 ( .A1(n586), .A2(n649), .ZN(n669) );
  INV_X1 U665 ( .A(n669), .ZN(n587) );
  NOR2_X1 U666 ( .A1(n720), .A2(n587), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT49), .B(n597), .Z(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n602), .B(KEYINPUT119), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U675 ( .A(n608), .B(KEYINPUT120), .ZN(n609) );
  NOR2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n614) );
  NOR2_X1 U677 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U679 ( .A1(n615), .A2(n621), .ZN(n616) );
  NOR2_X1 U680 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U681 ( .A(n618), .B(KEYINPUT52), .ZN(n620) );
  NOR2_X1 U682 ( .A1(n620), .A2(n619), .ZN(n624) );
  NOR2_X1 U683 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U684 ( .A(KEYINPUT53), .B(n626), .Z(G75) );
  NAND2_X1 U685 ( .A1(n670), .A2(G472), .ZN(n631) );
  XOR2_X1 U686 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n628) );
  XNOR2_X1 U687 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U688 ( .A(n631), .B(n630), .ZN(n634) );
  INV_X1 U689 ( .A(G952), .ZN(n632) );
  NAND2_X1 U690 ( .A1(n632), .A2(G953), .ZN(n633) );
  NAND2_X1 U691 ( .A1(n634), .A2(n676), .ZN(n635) );
  XNOR2_X1 U692 ( .A(n635), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U693 ( .A1(n670), .A2(G475), .ZN(n639) );
  XNOR2_X1 U694 ( .A(KEYINPUT87), .B(KEYINPUT59), .ZN(n636) );
  XNOR2_X1 U695 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U696 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U697 ( .A1(n640), .A2(n676), .ZN(n642) );
  XOR2_X1 U698 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n641) );
  XNOR2_X1 U699 ( .A(n642), .B(n641), .ZN(G60) );
  BUF_X2 U700 ( .A(n670), .Z(n687) );
  NAND2_X1 U701 ( .A1(n687), .A2(G478), .ZN(n645) );
  XNOR2_X1 U702 ( .A(n643), .B(KEYINPUT125), .ZN(n644) );
  XNOR2_X1 U703 ( .A(n645), .B(n644), .ZN(n646) );
  INV_X1 U704 ( .A(n676), .ZN(n691) );
  NOR2_X1 U705 ( .A1(n646), .A2(n691), .ZN(G63) );
  XNOR2_X1 U706 ( .A(KEYINPUT114), .B(n647), .ZN(G3) );
  NOR2_X1 U707 ( .A1(n650), .A2(n661), .ZN(n648) );
  XOR2_X1 U708 ( .A(G104), .B(n648), .Z(G6) );
  INV_X1 U709 ( .A(n649), .ZN(n664) );
  NOR2_X1 U710 ( .A1(n650), .A2(n664), .ZN(n652) );
  XNOR2_X1 U711 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n651) );
  XNOR2_X1 U712 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U713 ( .A(n344), .B(n653), .ZN(G9) );
  XOR2_X1 U714 ( .A(G110), .B(n654), .Z(G12) );
  NOR2_X1 U715 ( .A1(n664), .A2(n658), .ZN(n656) );
  XNOR2_X1 U716 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n655) );
  XNOR2_X1 U717 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U718 ( .A(G128), .B(n657), .Z(G30) );
  NOR2_X1 U719 ( .A1(n661), .A2(n658), .ZN(n659) );
  XOR2_X1 U720 ( .A(KEYINPUT116), .B(n659), .Z(n660) );
  XNOR2_X1 U721 ( .A(G146), .B(n660), .ZN(G48) );
  NOR2_X1 U722 ( .A1(n661), .A2(n663), .ZN(n662) );
  XOR2_X1 U723 ( .A(G113), .B(n662), .Z(G15) );
  NOR2_X1 U724 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U725 ( .A(G116), .B(n665), .Z(G18) );
  XOR2_X1 U726 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n668) );
  XNOR2_X1 U727 ( .A(n666), .B(G125), .ZN(n667) );
  XNOR2_X1 U728 ( .A(n668), .B(n667), .ZN(G27) );
  XNOR2_X1 U729 ( .A(G134), .B(n669), .ZN(G36) );
  NAND2_X1 U730 ( .A1(n670), .A2(G210), .ZN(n675) );
  XOR2_X1 U731 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n673) );
  XNOR2_X1 U732 ( .A(n671), .B(KEYINPUT85), .ZN(n672) );
  XNOR2_X1 U733 ( .A(n675), .B(n674), .ZN(n677) );
  NAND2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n680) );
  XOR2_X1 U735 ( .A(KEYINPUT80), .B(KEYINPUT122), .Z(n678) );
  XNOR2_X1 U736 ( .A(KEYINPUT56), .B(n678), .ZN(n679) );
  XNOR2_X1 U737 ( .A(n680), .B(n679), .ZN(G51) );
  NAND2_X1 U738 ( .A1(n687), .A2(G469), .ZN(n685) );
  XOR2_X1 U739 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  XNOR2_X1 U740 ( .A(n681), .B(KEYINPUT123), .ZN(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U743 ( .A1(n691), .A2(n686), .ZN(G54) );
  NAND2_X1 U744 ( .A1(n687), .A2(G217), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n692), .B(G101), .ZN(n693) );
  NAND2_X1 U746 ( .A1(n695), .A2(n694), .ZN(n703) );
  NOR2_X1 U747 ( .A1(n696), .A2(G953), .ZN(n701) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n697) );
  XOR2_X1 U749 ( .A(KEYINPUT61), .B(n697), .Z(n698) );
  NOR2_X1 U750 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U751 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U753 ( .A(KEYINPUT126), .B(n704), .ZN(G69) );
  XOR2_X1 U754 ( .A(n706), .B(n705), .Z(n707) );
  XNOR2_X1 U755 ( .A(n708), .B(n707), .ZN(n712) );
  XNOR2_X1 U756 ( .A(n712), .B(n709), .ZN(n711) );
  NAND2_X1 U757 ( .A1(n711), .A2(n710), .ZN(n716) );
  XNOR2_X1 U758 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U759 ( .A1(n713), .A2(G900), .ZN(n714) );
  NAND2_X1 U760 ( .A1(n714), .A2(G953), .ZN(n715) );
  NAND2_X1 U761 ( .A1(n716), .A2(n715), .ZN(G72) );
  XOR2_X1 U762 ( .A(G143), .B(n717), .Z(G45) );
  XOR2_X1 U763 ( .A(G137), .B(n718), .Z(G39) );
  XOR2_X1 U764 ( .A(n719), .B(G131), .Z(G33) );
  XOR2_X1 U765 ( .A(G140), .B(n720), .Z(G42) );
  XNOR2_X1 U766 ( .A(G119), .B(n721), .ZN(G21) );
endmodule

