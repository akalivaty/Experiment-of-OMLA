//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT2), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT80), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(new_n208), .A3(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n207), .B1(new_n215), .B2(KEYINPUT81), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n210), .A2(new_n212), .A3(new_n217), .A4(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(new_n214), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n209), .A2(new_n214), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(new_n204), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n205), .A2(new_n206), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n216), .A2(new_n218), .B1(new_n224), .B2(new_n225), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT82), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT76), .B(G218gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT22), .B1(new_n233), .B2(G211gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G197gat), .B(G204gat), .Z(new_n237));
  OR3_X1    g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n234), .B2(new_n237), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT87), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT87), .A4(new_n243), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n232), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n227), .B2(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G228gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n238), .A2(new_n240), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n258), .A2(new_n249), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n227), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n255), .B1(new_n260), .B2(new_n252), .ZN(new_n261));
  OAI21_X1  g060(.A(G22gat), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263));
  INV_X1    g062(.A(new_n261), .ZN(new_n264));
  INV_X1    g063(.A(G22gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n264), .B(new_n265), .C1(new_n248), .C2(new_n256), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT31), .B(G50gat), .Z(new_n268));
  XNOR2_X1  g067(.A(G78gat), .B(G106gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n267), .A2(new_n271), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(new_n266), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT88), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n229), .A2(new_n231), .A3(new_n277), .A4(KEYINPUT3), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G134gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n283), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(KEYINPUT1), .B2(new_n279), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n219), .A2(new_n226), .A3(KEYINPUT82), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT82), .B1(new_n219), .B2(new_n226), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT83), .B1(new_n230), .B2(new_n292), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n278), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n283), .A2(new_n282), .A3(new_n285), .ZN(new_n296));
  XOR2_X1   g095(.A(G113gat), .B(G120gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n282), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n296), .A2(new_n281), .B1(new_n298), .B2(new_n287), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n289), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n303), .A2(new_n304), .A3(new_n227), .ZN(new_n305));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT4), .B1(new_n230), .B2(new_n299), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n295), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n229), .A2(new_n231), .A3(new_n289), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n219), .A2(new_n226), .A3(new_n299), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n314), .B2(new_n307), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n302), .A3(new_n230), .A4(new_n304), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT85), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n323), .A2(new_n295), .A3(new_n306), .A4(new_n311), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G1gat), .B(G29gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT0), .ZN(new_n327));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT6), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n329), .A3(new_n324), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT38), .ZN(new_n335));
  OR3_X1    g134(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n342), .A2(KEYINPUT28), .A3(new_n341), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n342), .B2(new_n341), .ZN(new_n344));
  OAI221_X1 g143(.A(new_n339), .B1(new_n340), .B2(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT24), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n340), .B2(new_n341), .ZN(new_n347));
  NAND3_X1  g146(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n347), .B(new_n348), .C1(G183gat), .C2(G190gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n337), .B(KEYINPUT67), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351));
  OR3_X1    g150(.A1(new_n351), .A2(G169gat), .A3(G176gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT25), .ZN(new_n355));
  NOR2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT65), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(KEYINPUT64), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT64), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n346), .C1(new_n340), .C2(new_n341), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n358), .A2(new_n348), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n353), .A2(new_n363), .A3(new_n337), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT66), .B(G169gat), .Z(new_n365));
  NOR2_X1   g164(.A1(new_n351), .A2(G176gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n355), .A3(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n369), .B2(new_n249), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n251), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n251), .ZN(new_n375));
  AOI22_X1  g174(.A1(KEYINPUT25), .A2(new_n354), .B1(new_n362), .B2(new_n367), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n376), .B2(new_n345), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n375), .B(new_n371), .C1(new_n377), .C2(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(KEYINPUT37), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(KEYINPUT37), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n335), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n374), .A2(new_n378), .A3(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n383), .B1(new_n379), .B2(KEYINPUT37), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n375), .B1(new_n372), .B2(new_n373), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n371), .B(new_n251), .C1(new_n377), .C2(new_n370), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(KEYINPUT37), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n335), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n389), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n329), .B1(new_n316), .B2(new_n324), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n397), .A2(KEYINPUT86), .A3(KEYINPUT6), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT86), .B1(new_n397), .B2(KEYINPUT6), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n334), .B(new_n396), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n389), .ZN(new_n401));
  OR3_X1    g200(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n383), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n397), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT39), .B1(new_n314), .B2(new_n307), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n306), .B1(new_n323), .B2(new_n295), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT39), .B(new_n306), .C1(new_n323), .C2(new_n295), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n330), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT89), .A3(new_n329), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n410), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT91), .B(KEYINPUT40), .Z(new_n418));
  OAI21_X1  g217(.A(new_n404), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT40), .ZN(new_n420));
  AOI211_X1 g219(.A(new_n420), .B(new_n410), .C1(new_n416), .C2(new_n413), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n276), .B(new_n400), .C1(new_n419), .C2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n334), .B1(new_n398), .B2(new_n399), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n403), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n275), .A2(new_n267), .A3(new_n271), .ZN(new_n425));
  INV_X1    g224(.A(new_n272), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n303), .A2(new_n369), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n345), .A2(new_n376), .B1(new_n300), .B2(new_n302), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT72), .ZN(new_n435));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT33), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(KEYINPUT32), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(KEYINPUT70), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT70), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n303), .A2(new_n369), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n376), .A2(new_n300), .A3(new_n302), .A4(new_n345), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n429), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(KEYINPUT33), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n448), .A3(KEYINPUT32), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT32), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT71), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n451), .A3(new_n437), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n439), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n429), .A3(new_n444), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT34), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n429), .B2(KEYINPUT74), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n454), .B(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n428), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n457), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n446), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n460), .A2(new_n437), .A3(new_n449), .A4(new_n451), .ZN(new_n461));
  INV_X1    g260(.A(new_n457), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(KEYINPUT75), .A3(new_n462), .A4(new_n439), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(KEYINPUT73), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n453), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n424), .A2(new_n427), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n425), .A3(new_n426), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n424), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n473), .A2(new_n403), .A3(new_n276), .A4(new_n423), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n422), .A2(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(G1gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT16), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(G1gat), .B2(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G8gat), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n479), .B(new_n482), .C1(G1gat), .C2(new_n476), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n485));
  INV_X1    g284(.A(G29gat), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G50gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G43gat), .ZN(new_n492));
  INV_X1    g291(.A(G43gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G50gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT15), .ZN(new_n495));
  NAND2_X1  g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT96), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(G29gat), .A3(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n490), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n493), .A2(KEYINPUT94), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G43gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n491), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(G50gat), .B1(new_n502), .B2(new_n504), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT95), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n501), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n489), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT93), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n488), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n495), .B1(new_n517), .B2(new_n496), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n484), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT97), .ZN(new_n523));
  AND4_X1   g322(.A1(new_n523), .A2(new_n513), .A3(KEYINPUT17), .A4(new_n519), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n507), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n518), .B1(new_n525), .B2(new_n501), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(KEYINPUT17), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n522), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n484), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n532), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n484), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n529), .B(KEYINPUT13), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT12), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n535), .A2(new_n536), .A3(new_n542), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT98), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n541), .B1(new_n533), .B2(new_n534), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n536), .A4(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n536), .ZN(new_n554));
  INV_X1    g353(.A(new_n548), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n550), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n475), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n331), .B2(new_n332), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n397), .A2(KEYINPUT86), .A3(KEYINPUT6), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n397), .A2(KEYINPUT6), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n559), .A2(new_n560), .B1(new_n333), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT7), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n520), .B2(new_n521), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n524), .B2(new_n527), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n520), .A2(new_n580), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n564), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT103), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT102), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n579), .B1(new_n526), .B2(KEYINPUT17), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT97), .B1(new_n520), .B2(new_n521), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n526), .A2(new_n523), .A3(KEYINPUT17), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n584), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n563), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n582), .A2(new_n564), .A3(new_n584), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(KEYINPUT103), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n587), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n587), .B2(new_n595), .ZN(new_n600));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n595), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n596), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n601), .B1(new_n605), .B2(new_n598), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608));
  INV_X1    g407(.A(G57gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G64gat), .ZN(new_n610));
  INV_X1    g409(.A(G64gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(G57gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G71gat), .B(G78gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n616), .B2(new_n613), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n608), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G71gat), .A2(G78gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G57gat), .B(G64gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(new_n615), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT99), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT21), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n530), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT101), .ZN(new_n636));
  INV_X1    g435(.A(new_n632), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n637), .A3(new_n630), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n633), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n633), .B2(new_n638), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G183gat), .B(G211gat), .Z(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n639), .B2(new_n640), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n619), .A2(new_n579), .A3(new_n626), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n624), .A2(new_n625), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n574), .A2(KEYINPUT104), .A3(new_n576), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n576), .A2(KEYINPUT104), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n651), .A2(new_n578), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n650), .A2(new_n654), .A3(KEYINPUT105), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n580), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n650), .A2(new_n654), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n667), .A3(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n607), .A2(new_n649), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n557), .A2(new_n562), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  INV_X1    g479(.A(new_n557), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  INV_X1    g481(.A(new_n403), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n482), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n681), .A2(new_n403), .A3(new_n677), .A4(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(KEYINPUT42), .B2(new_n686), .ZN(G1325gat));
  INV_X1    g487(.A(new_n464), .ZN(new_n689));
  AOI21_X1  g488(.A(G15gat), .B1(new_n682), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n466), .A2(new_n469), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT106), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n690), .B1(new_n682), .B2(new_n694), .ZN(G1326gat));
  NAND3_X1  g494(.A1(new_n557), .A2(new_n427), .A3(new_n678), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n472), .A2(new_n474), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n427), .B1(new_n562), .B2(new_n683), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n422), .A2(new_n701), .A3(new_n691), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n550), .A2(new_n553), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n554), .A2(new_n555), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n607), .A2(new_n649), .A3(new_n675), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n486), .A3(new_n562), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n603), .A2(new_n606), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n703), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g515(.A(new_n607), .B(new_n712), .C1(new_n700), .C2(new_n702), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n649), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n675), .B(KEYINPUT108), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n706), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT109), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n718), .A2(new_n423), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n710), .B1(new_n724), .B2(new_n486), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n487), .A3(new_n683), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT46), .Z(new_n727));
  NOR3_X1   g526(.A1(new_n718), .A2(new_n403), .A3(new_n723), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n487), .B2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(new_n714), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n475), .B2(new_n607), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n703), .A2(new_n715), .A3(new_n711), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n733), .A2(new_n692), .B1(new_n502), .B2(new_n504), .ZN(new_n734));
  INV_X1    g533(.A(new_n708), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n464), .A3(new_n505), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n734), .B2(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n491), .B1(new_n733), .B2(new_n427), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n276), .A2(G50gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n708), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n427), .B(new_n722), .C1(new_n716), .C2(new_n717), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(KEYINPUT112), .A3(KEYINPUT48), .A4(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n747), .A2(new_n751), .A3(G50gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n747), .B2(G50gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n744), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n755), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g555(.A1(new_n715), .A2(new_n719), .A3(new_n720), .A4(new_n706), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n703), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n423), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n609), .ZN(G1332gat));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n403), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  OAI21_X1  g564(.A(KEYINPUT113), .B1(new_n758), .B2(new_n464), .ZN(new_n766));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n758), .A2(KEYINPUT113), .A3(new_n464), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n692), .A2(G71gat), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n768), .A2(new_n769), .B1(new_n758), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g571(.A1(new_n758), .A2(new_n276), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g573(.A1(new_n475), .A2(new_n607), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n649), .A2(new_n706), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n562), .A2(new_n571), .A3(new_n675), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n776), .A2(new_n675), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n718), .A2(new_n423), .A3(new_n784), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n782), .A2(new_n783), .B1(new_n785), .B2(new_n571), .ZN(G1336gat));
  NOR2_X1   g585(.A1(new_n403), .A2(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n720), .B(new_n788), .C1(new_n779), .C2(new_n780), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n718), .A2(new_n784), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n572), .B1(new_n790), .B2(new_n683), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT52), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n720), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n781), .A2(new_n793), .A3(new_n787), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n718), .A2(new_n403), .A3(new_n784), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n794), .B(new_n795), .C1(new_n572), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n797), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n689), .A2(new_n799), .A3(new_n675), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n718), .A2(new_n691), .A3(new_n784), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n782), .A2(new_n800), .B1(new_n801), .B2(new_n799), .ZN(G1338gat));
  NOR2_X1   g601(.A1(new_n276), .A2(G106gat), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n720), .B(new_n804), .C1(new_n779), .C2(new_n780), .ZN(new_n805));
  INV_X1    g604(.A(G106gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n790), .B2(new_n427), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT53), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n781), .A2(new_n793), .A3(new_n803), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n718), .A2(new_n276), .A3(new_n784), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n809), .B(new_n810), .C1(new_n806), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n660), .A2(new_n666), .A3(new_n661), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n661), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n658), .B2(new_n659), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n666), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n816), .A2(new_n664), .A3(KEYINPUT54), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n666), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n671), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n674), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n827), .A3(new_n674), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n666), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT54), .B1(new_n818), .B2(new_n666), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT114), .B1(new_n818), .B2(new_n666), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n672), .B1(new_n664), .B2(KEYINPUT54), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n826), .A2(new_n706), .A3(new_n828), .A4(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n531), .A2(new_n537), .A3(new_n539), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT116), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n528), .A2(new_n532), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n529), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n547), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n704), .A2(new_n675), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n715), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n550), .A2(new_n553), .B1(new_n840), .B2(new_n547), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n603), .B2(new_n606), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n827), .B1(new_n824), .B2(new_n674), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n835), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n719), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n677), .A2(new_n706), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n423), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n471), .A2(new_n683), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n706), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n427), .B1(new_n849), .B2(new_n851), .ZN(new_n857));
  AND4_X1   g656(.A1(new_n403), .A2(new_n857), .A3(new_n562), .A4(new_n689), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n706), .A2(G113gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  NAND3_X1  g659(.A1(new_n858), .A2(G120gat), .A3(new_n793), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n284), .B1(new_n854), .B2(new_n676), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT117), .ZN(G1341gat));
  NAND3_X1  g663(.A1(new_n858), .A2(G127gat), .A3(new_n649), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  AOI21_X1  g667(.A(G127gat), .B1(new_n855), .B2(new_n649), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1342gat));
  OR3_X1    g669(.A1(new_n854), .A2(G134gat), .A3(new_n607), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n858), .A2(new_n715), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G134gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n692), .A2(new_n683), .A3(new_n423), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n847), .A2(new_n846), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n715), .A3(new_n844), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n835), .A2(new_n674), .A3(new_n824), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT120), .B(new_n842), .C1(new_n880), .C2(new_n556), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n607), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n706), .A2(new_n674), .A3(new_n824), .A4(new_n835), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT120), .B1(new_n883), .B2(new_n842), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n850), .B1(new_n885), .B2(new_n719), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n276), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n849), .A2(new_n851), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n427), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n706), .B(new_n877), .C1(new_n888), .C2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT122), .B1(new_n893), .B2(G141gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n276), .B1(new_n466), .B2(new_n469), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n403), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n896), .B2(new_n895), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n208), .A2(new_n898), .A3(new_n706), .A4(new_n852), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n893), .B2(G141gat), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n894), .A2(new_n900), .A3(KEYINPUT58), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  AOI221_X4 g701(.A(new_n899), .B1(KEYINPUT122), .B2(new_n902), .C1(new_n893), .C2(G141gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(G1344gat));
  XOR2_X1   g703(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n905));
  NAND2_X1  g704(.A1(new_n877), .A2(new_n675), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n886), .A2(new_n276), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n887), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n276), .B1(new_n849), .B2(new_n851), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n890), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n905), .B1(new_n911), .B2(new_n213), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n675), .B(new_n877), .C1(new_n888), .C2(new_n892), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n213), .A2(KEYINPUT59), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(KEYINPUT123), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT123), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n898), .A2(new_n852), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n213), .A3(new_n675), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(new_n877), .B1(new_n888), .B2(new_n892), .ZN(new_n921));
  OAI21_X1  g720(.A(G155gat), .B1(new_n921), .B2(new_n719), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n202), .A3(new_n649), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n921), .B2(new_n607), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n918), .A2(new_n203), .A3(new_n715), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n562), .A2(new_n403), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n464), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n857), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n556), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n562), .B1(new_n849), .B2(new_n851), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n471), .A2(new_n403), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n706), .A2(new_n365), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n931), .B2(new_n720), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n676), .A2(G176gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n935), .B2(new_n939), .ZN(G1349gat));
  OAI21_X1  g739(.A(G183gat), .B1(new_n931), .B2(new_n719), .ZN(new_n941));
  INV_X1    g740(.A(new_n935), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n649), .A2(new_n342), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n942), .A2(KEYINPUT125), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT125), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n341), .A3(new_n715), .ZN(new_n949));
  OAI21_X1  g748(.A(G190gat), .B1(new_n931), .B2(new_n607), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1351gat));
  AND3_X1   g752(.A1(new_n933), .A2(new_n683), .A3(new_n895), .ZN(new_n954));
  XNOR2_X1  g753(.A(KEYINPUT126), .B(G197gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n706), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n907), .A2(new_n887), .B1(new_n909), .B2(new_n890), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n692), .A2(new_n929), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n957), .A2(new_n556), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n960), .B2(new_n955), .ZN(G1352gat));
  INV_X1    g760(.A(G204gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n954), .A2(new_n962), .A3(new_n675), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT62), .Z(new_n964));
  NOR3_X1   g763(.A1(new_n957), .A2(new_n720), .A3(new_n959), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR4_X1   g766(.A1(new_n957), .A2(KEYINPUT127), .A3(new_n720), .A4(new_n959), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1353gat));
  INV_X1    g768(.A(G211gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n970), .A3(new_n649), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n886), .A2(new_n276), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(KEYINPUT57), .ZN(new_n973));
  INV_X1    g772(.A(new_n910), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n649), .B(new_n958), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  AOI21_X1  g777(.A(G218gat), .B1(new_n954), .B2(new_n715), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n957), .A2(new_n959), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n715), .A2(new_n233), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(G1355gat));
endmodule


