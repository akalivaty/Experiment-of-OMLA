//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1151, new_n1152, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1219, new_n1220;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G97), .A2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G226), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n202), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G58), .A2(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n208), .B(new_n214), .C1(G107), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT66), .B(G77), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n232), .A2(G50), .A3(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n224), .B(new_n228), .C1(new_n231), .C2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n213), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  INV_X1    g0047(.A(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n212), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n229), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT7), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G20), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n216), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G58), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n216), .ZN(new_n268));
  OAI21_X1  g0068(.A(G20), .B1(new_n268), .B2(new_n201), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G159), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n266), .A2(KEYINPUT16), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT7), .B1(new_n263), .B2(new_n264), .ZN(new_n275));
  NOR4_X1   g0075(.A1(new_n261), .A2(new_n262), .A3(new_n258), .A4(G20), .ZN(new_n276));
  OAI21_X1  g0076(.A(G68), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n272), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n257), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n282), .A2(new_n264), .A3(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n257), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G1), .B2(new_n264), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n286), .B2(new_n281), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  INV_X1    g0089(.A(G1), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT69), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G1698), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n259), .A3(G223), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G87), .ZN(new_n300));
  OAI211_X1 g0100(.A(G226), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G33), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  OAI211_X1 g0104(.A(G1), .B(G13), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n293), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n291), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G232), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n280), .A2(new_n288), .B1(new_n289), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n302), .A2(new_n306), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  INV_X1    g0114(.A(new_n293), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n310), .A4(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n307), .A2(KEYINPUT75), .A3(new_n314), .A4(new_n310), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT18), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n311), .A2(G200), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n307), .A2(G190), .A3(new_n310), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n280), .A2(new_n323), .A3(new_n324), .A4(new_n288), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT17), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n283), .A2(new_n202), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n264), .A2(G33), .ZN(new_n330));
  INV_X1    g0130(.A(G150), .ZN(new_n331));
  INV_X1    g0131(.A(new_n270), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n281), .A2(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G20), .B2(new_n203), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n329), .B1(new_n202), .B2(new_n286), .C1(new_n334), .C2(new_n285), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G223), .A2(G1698), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT69), .B(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(G222), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n259), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n306), .C1(new_n219), .C2(new_n259), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n315), .C1(new_n207), .C2(new_n308), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n335), .A2(new_n336), .B1(G200), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT10), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n335), .B1(new_n343), .B2(G179), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n343), .A2(new_n289), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n263), .A2(new_n294), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G238), .B1(G107), .B2(new_n263), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n298), .A2(new_n259), .A3(G232), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n306), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n309), .A2(G244), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n357), .A2(new_n314), .A3(new_n315), .A4(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n286), .A2(new_n253), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n219), .A2(G20), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n361), .B1(new_n332), .B2(new_n281), .C1(new_n330), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(new_n257), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n220), .A2(new_n283), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n357), .A2(new_n315), .A3(new_n358), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n289), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(G200), .ZN(new_n371));
  INV_X1    g0171(.A(new_n366), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n372), .C1(new_n345), .C2(new_n368), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n348), .A2(new_n352), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT70), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n375), .A2(new_n376), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n303), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n295), .A2(new_n297), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT71), .B1(new_n387), .B2(G226), .ZN(new_n388));
  AND4_X1   g0188(.A1(KEYINPUT71), .A2(new_n298), .A3(new_n259), .A4(G226), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n382), .B(new_n383), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n306), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n293), .B(KEYINPUT72), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n305), .B2(new_n291), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n393), .A2(new_n217), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AND4_X1   g0197(.A1(new_n381), .A2(new_n391), .A3(new_n392), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n390), .B2(new_n306), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n381), .B1(new_n399), .B2(new_n392), .ZN(new_n400));
  OAI211_X1 g0200(.A(G169), .B(new_n380), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n391), .A2(new_n392), .A3(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT13), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n381), .A3(new_n392), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(G179), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n289), .B1(new_n403), .B2(new_n404), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n401), .B(new_n405), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n216), .A2(G20), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n409), .B1(new_n330), .B2(new_n253), .C1(new_n332), .C2(new_n202), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n216), .B2(new_n286), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n283), .A2(new_n216), .ZN(new_n413));
  XOR2_X1   g0213(.A(new_n413), .B(KEYINPUT12), .Z(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT11), .B1(new_n410), .B2(new_n257), .ZN(new_n415));
  OR3_X1    g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n398), .A2(new_n400), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G190), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n403), .A2(new_n404), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(G200), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n408), .A2(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AND4_X1   g0221(.A1(new_n328), .A2(new_n377), .A3(new_n378), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G116), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n353), .A2(G244), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT77), .B1(new_n387), .B2(G238), .ZN(new_n425));
  AND4_X1   g0225(.A1(KEYINPUT77), .A2(new_n298), .A3(new_n259), .A4(G238), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n306), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n290), .A2(G45), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n292), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n305), .A2(G250), .A3(new_n429), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n428), .A2(new_n314), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n259), .A2(new_n264), .A3(G68), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT19), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n264), .B1(new_n382), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(G97), .A2(G107), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n210), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n382), .B2(G20), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n434), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n257), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n362), .A2(new_n283), .ZN(new_n443));
  INV_X1    g0243(.A(new_n283), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n285), .C1(G1), .C2(new_n303), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(new_n443), .C1(new_n362), .C2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n432), .ZN(new_n447));
  AOI211_X1 g0247(.A(new_n430), .B(new_n447), .C1(new_n427), .C2(new_n306), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n433), .B(new_n446), .C1(new_n448), .C2(G169), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n428), .A2(G190), .A3(new_n431), .A4(new_n432), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n445), .A2(new_n210), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n442), .A2(new_n443), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G200), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n450), .B(new_n452), .C1(new_n448), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT24), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(G20), .B2(new_n248), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT79), .B1(new_n423), .B2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(new_n264), .A3(G33), .A4(G116), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n456), .A2(new_n248), .A3(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n456), .A2(new_n248), .A3(KEYINPUT80), .A4(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT81), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n264), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT22), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n455), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT81), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT81), .B1(new_n461), .B2(new_n466), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n455), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n257), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n445), .A2(new_n248), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n444), .A2(G107), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n298), .A2(new_n259), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n211), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n306), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n290), .B(G45), .C1(new_n304), .C2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G41), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n305), .B(G264), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  OR3_X1    g0295(.A1(new_n493), .A2(KEYINPUT76), .A3(G41), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT76), .B1(new_n493), .B2(G41), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(G274), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n492), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n491), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n345), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n479), .A2(new_n481), .A3(new_n486), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n501), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n453), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n449), .B(new_n454), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT24), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n285), .B1(new_n509), .B2(new_n477), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n480), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n501), .A2(new_n314), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n499), .B1(new_n490), .B2(new_n306), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n289), .B1(new_n513), .B2(new_n495), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(KEYINPUT83), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n511), .A2(new_n486), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n283), .A2(new_n212), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  INV_X1    g0319(.A(G97), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n264), .C1(G33), .C2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n257), .C1(new_n264), .C2(G116), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT20), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  OAI221_X1 g0325(.A(new_n518), .B1(new_n212), .B2(new_n445), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n305), .B(G270), .C1(new_n492), .C2(new_n494), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT78), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n259), .A2(new_n532), .A3(G264), .A4(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n298), .A2(new_n259), .A3(G257), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n263), .A2(G303), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n529), .B1(new_n536), .B2(new_n306), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(G190), .A3(new_n500), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n500), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n527), .B(new_n538), .C1(new_n540), .C2(new_n453), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(G179), .A3(new_n526), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n289), .B1(new_n537), .B2(new_n500), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(new_n526), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n543), .B2(new_n526), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n541), .B(new_n542), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n444), .A2(G97), .ZN(new_n548));
  OAI21_X1  g0348(.A(G107), .B1(new_n275), .B2(new_n276), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT6), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n520), .A2(new_n248), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n437), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n248), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n270), .A2(G77), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n549), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n548), .B1(new_n557), .B2(new_n257), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n520), .B2(new_n445), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n489), .B2(new_n218), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n387), .A2(KEYINPUT4), .A3(G244), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n353), .A2(G250), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n519), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n306), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n305), .B(G257), .C1(new_n492), .C2(new_n494), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n565), .A2(new_n314), .A3(new_n500), .A4(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n566), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n499), .B(new_n568), .C1(new_n564), .C2(new_n306), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n559), .B(new_n567), .C1(new_n569), .C2(G169), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n445), .A2(new_n520), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n548), .B(new_n571), .C1(new_n557), .C2(new_n257), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(G190), .A3(new_n500), .A4(new_n566), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n569), .C2(new_n453), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR4_X1   g0375(.A1(new_n507), .A2(new_n517), .A3(new_n547), .A4(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n422), .A2(new_n576), .ZN(G372));
  NAND2_X1  g0377(.A1(new_n449), .A2(new_n454), .ZN(new_n578));
  INV_X1    g0378(.A(new_n506), .ZN(new_n579));
  NOR4_X1   g0379(.A1(new_n510), .A2(new_n480), .A3(new_n502), .A4(new_n485), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n570), .A2(new_n574), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n582), .C1(new_n517), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n449), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n449), .A2(new_n454), .ZN(new_n586));
  INV_X1    g0386(.A(new_n570), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(KEYINPUT26), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT26), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n578), .B2(new_n570), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n585), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n422), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n420), .A2(new_n418), .ZN(new_n594));
  INV_X1    g0394(.A(new_n416), .ZN(new_n595));
  OAI21_X1  g0395(.A(G169), .B1(new_n398), .B2(new_n400), .ZN(new_n596));
  INV_X1    g0396(.A(new_n407), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n417), .B2(G179), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n598), .B2(new_n401), .ZN(new_n599));
  INV_X1    g0399(.A(new_n370), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n326), .B(new_n594), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT18), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT84), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n312), .B2(new_n320), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n311), .A2(new_n289), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT16), .B1(new_n266), .B2(new_n272), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n277), .A2(new_n274), .A3(new_n278), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n285), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n287), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n318), .A2(new_n319), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT84), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n602), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n312), .A2(new_n320), .A3(new_n603), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT84), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT18), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n601), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n351), .B1(new_n617), .B2(new_n348), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n593), .A2(new_n618), .ZN(G369));
  AOI21_X1  g0419(.A(new_n517), .B1(new_n579), .B2(new_n580), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n511), .A2(new_n486), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n282), .A2(G20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n290), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT85), .Z(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(G213), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n620), .A2(new_n630), .B1(new_n517), .B2(new_n629), .ZN(new_n631));
  INV_X1    g0431(.A(new_n629), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n583), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n547), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n629), .A2(new_n526), .ZN(new_n636));
  MUX2_X1   g0436(.A(new_n583), .B(new_n635), .S(new_n636), .Z(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(G330), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n620), .A2(new_n583), .A3(new_n632), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n517), .A2(new_n632), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(G399));
  NOR2_X1   g0443(.A1(new_n438), .A2(G116), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n225), .A2(new_n304), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G1), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n234), .B2(new_n645), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT28), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n569), .A2(new_n505), .A3(G179), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n539), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n565), .A2(new_n500), .A3(new_n566), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n537), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n448), .A2(new_n569), .A3(new_n512), .A4(new_n537), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT30), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT31), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(new_n659), .A3(new_n629), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n658), .B2(new_n629), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT86), .ZN(new_n663));
  INV_X1    g0463(.A(new_n517), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n581), .A2(new_n664), .A3(new_n635), .A4(new_n582), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(new_n629), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n632), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n629), .B1(new_n584), .B2(new_n591), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT29), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(KEYINPUT87), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n670), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n648), .B1(new_n676), .B2(G1), .ZN(G364));
  NAND2_X1  g0477(.A1(new_n622), .A2(G45), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n645), .A2(G1), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT88), .Z(new_n680));
  NOR2_X1   g0480(.A1(new_n264), .A2(new_n314), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(G190), .A3(new_n453), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT89), .Z(new_n683));
  INV_X1    g0483(.A(new_n681), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n684), .A2(G190), .A3(G200), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n683), .A2(G58), .B1(new_n219), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(G190), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n453), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n202), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT90), .ZN(new_n691));
  NOR2_X1   g0491(.A1(G179), .A2(G200), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G190), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G20), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n693), .ZN(new_n697));
  INV_X1    g0497(.A(G159), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT32), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n264), .A2(G179), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n345), .A3(G200), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n248), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(G190), .A3(G200), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n684), .A2(new_n453), .A3(G190), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n259), .B1(new_n210), .B2(new_n706), .C1(new_n708), .C2(new_n216), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n701), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n699), .A2(new_n700), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n695), .A2(G97), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n691), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n685), .A2(G311), .B1(new_n688), .B2(G326), .ZN(new_n714));
  XOR2_X1   g0514(.A(KEYINPUT33), .B(G317), .Z(new_n715));
  INV_X1    g0515(.A(G283), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n714), .B1(new_n708), .B2(new_n715), .C1(new_n716), .C2(new_n704), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(G294), .B2(new_n695), .ZN(new_n718));
  INV_X1    g0518(.A(new_n697), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G329), .ZN(new_n720));
  INV_X1    g0520(.A(new_n682), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G322), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G303), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n263), .B1(new_n706), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT93), .Z(new_n726));
  OAI21_X1  g0526(.A(new_n713), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n229), .B1(G20), .B2(new_n289), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n680), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n729), .B1(new_n637), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n732), .A2(new_n728), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n263), .A2(new_n225), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n234), .A2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(G45), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n737), .B(new_n738), .C1(new_n254), .C2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n259), .A2(new_n225), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n740), .B1(G116), .B2(new_n225), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n734), .B1(new_n735), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n637), .A2(G330), .ZN(new_n746));
  INV_X1    g0546(.A(new_n638), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n680), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(G396));
  INV_X1    g0549(.A(KEYINPUT97), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n370), .B2(new_n632), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n367), .A2(KEYINPUT97), .A3(new_n369), .A4(new_n629), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n370), .B(new_n373), .C1(new_n372), .C2(new_n632), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT98), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT98), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n753), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n671), .B(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(new_n670), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n680), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n704), .A2(new_n210), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n719), .B2(G311), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n708), .A2(new_n716), .B1(new_n689), .B2(new_n724), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G116), .B2(new_n685), .ZN(new_n767));
  INV_X1    g0567(.A(new_n706), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n259), .B1(new_n768), .B2(G107), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n767), .A2(new_n712), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n765), .B(new_n770), .C1(new_n771), .C2(new_n682), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n683), .A2(G143), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G150), .A2(new_n707), .B1(new_n688), .B2(G137), .ZN(new_n774));
  INV_X1    g0574(.A(new_n685), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n773), .B(new_n774), .C1(new_n698), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT34), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n704), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G68), .B1(new_n695), .B2(G58), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n263), .B1(new_n768), .B2(G50), .ZN(new_n781));
  INV_X1    g0581(.A(G132), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n780), .B(new_n781), .C1(new_n782), .C2(new_n697), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT96), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT96), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n776), .A2(new_n777), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n772), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n680), .B1(new_n788), .B2(new_n728), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n728), .A2(new_n730), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(G77), .B2(new_n791), .C1(new_n759), .C2(new_n731), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n762), .A2(new_n792), .ZN(G384));
  AOI21_X1  g0593(.A(KEYINPUT86), .B1(new_n576), .B2(new_n632), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n511), .A2(new_n486), .A3(new_n579), .A4(new_n503), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n635), .A2(new_n582), .A3(new_n586), .A4(new_n795), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n796), .A2(new_n663), .A3(new_n517), .A4(new_n629), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n794), .A2(new_n797), .B1(new_n661), .B2(new_n660), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n408), .A2(new_n416), .A3(new_n629), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT100), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n629), .A2(new_n416), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n421), .A2(new_n802), .B1(new_n599), .B2(new_n629), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n803), .B2(new_n800), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT38), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n280), .A2(new_n288), .ZN(new_n806));
  INV_X1    g0606(.A(new_n627), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n321), .B(new_n602), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n326), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n321), .A2(new_n325), .A3(new_n808), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT37), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n805), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n811), .B(KEYINPUT37), .ZN(new_n815));
  OAI211_X1 g0615(.A(KEYINPUT38), .B(new_n815), .C1(new_n328), .C2(new_n808), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n798), .A2(new_n804), .A3(new_n759), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT40), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n759), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n408), .A2(new_n416), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n594), .A3(new_n802), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n800), .B1(new_n823), .B2(new_n799), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n821), .B1(new_n825), .B2(new_n801), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n808), .B1(new_n616), .B2(new_n326), .ZN(new_n827));
  INV_X1    g0627(.A(new_n325), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n613), .B2(new_n614), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT101), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n808), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(KEYINPUT101), .B(new_n828), .C1(new_n613), .C2(new_n614), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT37), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n811), .A2(KEYINPUT37), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n827), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n816), .B1(new_n835), .B2(KEYINPUT38), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n826), .A2(new_n836), .A3(KEYINPUT40), .A4(new_n798), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n820), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n422), .A2(new_n798), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G330), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT39), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n816), .C1(new_n835), .C2(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n822), .A2(new_n629), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n843), .A2(new_n848), .A3(new_n844), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n612), .A2(new_n615), .A3(new_n627), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n671), .A2(new_n759), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n370), .B2(new_n629), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n817), .A3(new_n804), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n841), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n422), .B1(new_n673), .B2(new_n675), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n618), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT103), .Z(new_n859));
  XNOR2_X1  g0659(.A(new_n856), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n290), .B2(new_n622), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n219), .B1(new_n267), .B2(new_n216), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n234), .A2(new_n862), .B1(G50), .B2(new_n216), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n282), .ZN(new_n864));
  OAI211_X1 g0664(.A(G20), .B(new_n230), .C1(new_n554), .C2(KEYINPUT35), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n212), .B(new_n865), .C1(KEYINPUT35), .C2(new_n554), .ZN(new_n866));
  XNOR2_X1  g0666(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n864), .A3(new_n868), .ZN(G367));
  NOR2_X1   g0669(.A1(new_n632), .A2(new_n452), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n585), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n578), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT43), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n587), .A2(new_n629), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n582), .B1(new_n572), .B2(new_n632), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n640), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT42), .Z(new_n877));
  OAI21_X1  g0677(.A(new_n570), .B1(new_n875), .B2(new_n664), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(new_n632), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n873), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n639), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n874), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n880), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n872), .A2(KEYINPUT43), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n884), .B(new_n885), .Z(new_n886));
  XNOR2_X1  g0686(.A(new_n645), .B(KEYINPUT41), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n639), .B(KEYINPUT105), .Z(new_n888));
  AOI21_X1  g0688(.A(new_n638), .B1(new_n634), .B2(new_n640), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n676), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n642), .A2(new_n882), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT104), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT45), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n893), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT45), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n642), .A2(new_n882), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT44), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n881), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n896), .A2(new_n899), .A3(new_n639), .A4(new_n901), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n892), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n887), .B1(new_n905), .B2(new_n676), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n678), .A2(G1), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n886), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n683), .A2(G303), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n695), .A2(G107), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n707), .A2(G294), .ZN(new_n911));
  INV_X1    g0711(.A(new_n703), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n688), .A2(G311), .B1(new_n912), .B2(G97), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n719), .A2(G317), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT46), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n706), .B2(new_n212), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n915), .A2(new_n263), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n914), .B(new_n919), .C1(G283), .C2(new_n685), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n688), .A2(G143), .ZN(new_n921));
  AOI22_X1  g0721(.A1(G50), .A2(new_n685), .B1(new_n707), .B2(G159), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT106), .Z(new_n923));
  AOI21_X1  g0723(.A(new_n263), .B1(new_n768), .B2(G58), .ZN(new_n924));
  AOI22_X1  g0724(.A1(G150), .A2(new_n721), .B1(new_n912), .B2(new_n219), .ZN(new_n925));
  INV_X1    g0725(.A(G137), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n924), .B(new_n925), .C1(new_n697), .C2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n696), .A2(new_n216), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n920), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT47), .Z(new_n931));
  AOI21_X1  g0731(.A(new_n680), .B1(new_n931), .B2(new_n728), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n735), .B1(new_n225), .B2(new_n362), .C1(new_n244), .C2(new_n736), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n932), .B(new_n933), .C1(new_n733), .C2(new_n872), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n908), .A2(new_n934), .ZN(G387));
  OAI22_X1  g0735(.A1(new_n696), .A2(new_n362), .B1(new_n520), .B2(new_n704), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n259), .B1(new_n220), .B2(new_n706), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n708), .A2(new_n281), .B1(new_n689), .B2(new_n698), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n682), .A2(new_n202), .ZN(new_n939));
  NOR4_X1   g0739(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(new_n216), .B2(new_n775), .C1(new_n331), .C2(new_n697), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n683), .A2(G317), .B1(G303), .B2(new_n685), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT111), .Z(new_n943));
  AOI22_X1  g0743(.A1(G311), .A2(new_n707), .B1(new_n688), .B2(G322), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT112), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT48), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n695), .A2(G283), .B1(G294), .B2(new_n768), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT110), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT49), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT49), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n259), .B1(new_n719), .B2(G326), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n703), .A2(new_n212), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n941), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n680), .B1(new_n956), .B2(new_n728), .ZN(new_n957));
  INV_X1    g0757(.A(new_n631), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n958), .B2(new_n733), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n281), .A2(G50), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n644), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  AOI21_X1  g0764(.A(G45), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n962), .B(new_n965), .C1(new_n964), .C2(new_n963), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n216), .A2(new_n253), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n737), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT109), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n739), .B2(new_n241), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(G107), .B2(new_n225), .C1(new_n644), .C2(new_n742), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n959), .B1(new_n735), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n890), .B2(new_n907), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n645), .B(KEYINPUT113), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n892), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n676), .B2(new_n890), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(G393));
  INV_X1    g0777(.A(new_n974), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n905), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n903), .A2(new_n904), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n892), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n907), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n263), .B1(new_n716), .B2(new_n706), .C1(new_n775), .C2(new_n771), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n705), .B(new_n983), .C1(new_n719), .C2(G322), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G317), .A2(new_n688), .B1(new_n721), .B2(G311), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n696), .A2(new_n212), .B1(new_n985), .B2(KEYINPUT52), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(KEYINPUT52), .B2(new_n985), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n984), .B(new_n987), .C1(new_n724), .C2(new_n708), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT114), .Z(new_n989));
  OAI221_X1 g0789(.A(new_n259), .B1(new_n708), .B2(new_n202), .C1(new_n281), .C2(new_n775), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n763), .B(new_n990), .C1(new_n719), .C2(G143), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G150), .A2(new_n688), .B1(new_n721), .B2(G159), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT51), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G77), .B2(new_n695), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n991), .B(new_n994), .C1(new_n216), .C2(new_n706), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n680), .B1(new_n996), .B2(new_n728), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n735), .B1(new_n520), .B2(new_n225), .C1(new_n250), .C2(new_n736), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(new_n733), .C2(new_n882), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n982), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n981), .A2(new_n1000), .ZN(G390));
  AND4_X1   g0801(.A1(G330), .A2(new_n798), .A3(new_n759), .A4(new_n804), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n847), .B1(new_n853), .B2(new_n804), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n846), .B2(new_n849), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n801), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT115), .B1(new_n824), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT115), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(new_n801), .C1(new_n803), .C2(new_n800), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n853), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n847), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n836), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1002), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n836), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1002), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n843), .A2(new_n848), .A3(new_n844), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n848), .B1(new_n843), .B2(new_n844), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1014), .B(new_n1015), .C1(new_n1018), .C2(new_n1003), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n422), .A2(G330), .A3(new_n798), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n857), .A2(new_n1021), .A3(new_n618), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n668), .A2(new_n669), .A3(new_n821), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT116), .B1(new_n1023), .B2(new_n1009), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n853), .B1(new_n670), .B2(new_n826), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n798), .A2(G330), .A3(new_n759), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT116), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n804), .B1(new_n670), .B2(new_n759), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n853), .B1(new_n1030), .B2(new_n1002), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1022), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1020), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1013), .A2(new_n1032), .A3(new_n1019), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n978), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(G125), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n259), .B1(new_n202), .B2(new_n703), .C1(new_n697), .C2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT117), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n768), .A2(G150), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT53), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n707), .A2(G137), .ZN(new_n1042));
  INV_X1    g0842(.A(G128), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT54), .B(G143), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1042), .B1(new_n689), .B2(new_n1043), .C1(new_n775), .C2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1041), .B(new_n1045), .C1(G159), .C2(new_n695), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1039), .B(new_n1046), .C1(new_n782), .C2(new_n682), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n696), .A2(new_n253), .B1(new_n216), .B2(new_n704), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n263), .B1(new_n706), .B2(new_n210), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n707), .A2(G107), .B1(new_n721), .B2(G116), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n520), .B2(new_n775), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n716), .B2(new_n689), .C1(new_n771), .C2(new_n697), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n680), .B1(new_n1054), .B2(new_n728), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1018), .B2(new_n731), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n281), .B2(new_n790), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1020), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n907), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1036), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT118), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1036), .A2(new_n1059), .A3(KEYINPUT118), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(G378));
  AND3_X1   g0864(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n820), .A2(new_n837), .A3(G330), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n807), .A2(new_n335), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n348), .A2(new_n352), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n348), .B2(new_n352), .ZN(new_n1069));
  OR3_X1    g0869(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT55), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT55), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1070), .A2(KEYINPUT56), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT56), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n820), .A2(new_n837), .A3(new_n1074), .A4(G330), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1065), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT120), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n855), .A2(new_n1077), .A3(new_n1076), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1065), .A2(new_n1078), .A3(KEYINPUT120), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n907), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n708), .A2(new_n782), .B1(new_n706), .B2(new_n1044), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n775), .A2(new_n926), .B1(new_n689), .B2(new_n1037), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G150), .C2(new_n695), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1043), .B2(new_n682), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT59), .Z(new_n1089));
  AOI21_X1  g0889(.A(G41), .B1(new_n719), .B2(G124), .ZN(new_n1090));
  AOI21_X1  g0890(.A(G33), .B1(new_n912), .B2(G159), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n263), .B1(new_n697), .B2(new_n716), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n362), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1094), .A2(new_n685), .B1(new_n707), .B2(G97), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n304), .C1(new_n220), .C2(new_n706), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n688), .A2(G116), .B1(new_n912), .B2(G58), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n248), .B2(new_n682), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1093), .A2(new_n928), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT58), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n261), .A2(G41), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1099), .A2(KEYINPUT58), .B1(G50), .B2(new_n1101), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1102), .A2(KEYINPUT119), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(KEYINPUT119), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1092), .A2(new_n1100), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n680), .B1(new_n1105), .B2(new_n728), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(G50), .B2(new_n791), .C1(new_n1075), .C2(new_n731), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1084), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1022), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1035), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1082), .A2(new_n1111), .A3(new_n1083), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT57), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT121), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1079), .A2(new_n1115), .A3(new_n1081), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1065), .A2(new_n1078), .A3(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1116), .A2(new_n1111), .A3(KEYINPUT57), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n978), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1109), .B1(new_n1114), .B2(new_n1119), .ZN(G375));
  NAND3_X1  g0920(.A1(new_n1029), .A2(new_n1031), .A3(new_n1022), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OR3_X1    g0922(.A1(new_n1122), .A2(new_n887), .A3(new_n1032), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n907), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n708), .A2(new_n1044), .B1(new_n698), .B2(new_n706), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G150), .B2(new_n685), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n683), .A2(G137), .B1(G50), .B2(new_n695), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n263), .B1(new_n912), .B2(G58), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n1043), .B2(new_n697), .C1(new_n782), .C2(new_n689), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n696), .A2(new_n362), .B1(new_n253), .B2(new_n704), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n263), .B1(new_n682), .B2(new_n716), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n708), .A2(new_n212), .B1(new_n520), .B2(new_n706), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n689), .A2(new_n771), .ZN(new_n1135));
  NOR4_X1   g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n248), .B2(new_n775), .C1(new_n724), .C2(new_n697), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT122), .Z(new_n1139));
  AOI21_X1  g0939(.A(new_n680), .B1(new_n1139), .B2(new_n728), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(G68), .B2(new_n791), .C1(new_n1009), .C2(new_n731), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT123), .B1(new_n1125), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1125), .A2(KEYINPUT123), .A3(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1123), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT124), .ZN(G381));
  NOR4_X1   g0945(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(G375), .A2(new_n1060), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n908), .A2(new_n934), .A3(new_n1000), .A4(new_n981), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(G407));
  INV_X1    g0950(.A(G213), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1147), .B2(new_n628), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(G407), .A2(new_n1152), .ZN(G409));
  NAND3_X1  g0953(.A1(new_n1116), .A2(new_n907), .A3(new_n1117), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1107), .B(new_n1154), .C1(new_n1112), .C2(new_n887), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1060), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1036), .A2(new_n1059), .A3(KEYINPUT118), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT118), .B1(new_n1036), .B2(new_n1059), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1157), .B1(G375), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT60), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n974), .B1(new_n1121), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1029), .A2(new_n1031), .A3(KEYINPUT60), .A4(new_n1022), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1033), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1166));
  INV_X1    g0966(.A(G384), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1165), .B(G384), .C1(new_n1143), .C2(new_n1142), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1151), .A2(G343), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1161), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT62), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT61), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT125), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT125), .ZN(new_n1178));
  INV_X1    g0978(.A(G2897), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1170), .A2(new_n1178), .B1(new_n1179), .B2(new_n1173), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1168), .A2(KEYINPUT125), .A3(new_n1169), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1177), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1118), .A2(new_n978), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1108), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1186), .A2(G378), .B1(new_n1156), .B2(new_n1155), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n1187), .B2(new_n1172), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT62), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1161), .A2(new_n1189), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1175), .A2(new_n1176), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(G387), .A2(G390), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(G393), .B(G396), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n1148), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1193), .B2(new_n1148), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1161), .A2(new_n1173), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT61), .B1(new_n1199), .B2(new_n1183), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT127), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n1175), .A3(new_n1201), .A4(new_n1190), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1192), .A2(new_n1198), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1183), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1185), .A2(new_n978), .A3(new_n1118), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(G378), .A2(new_n1205), .A3(new_n1109), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1172), .B1(new_n1206), .B2(new_n1157), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT63), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT61), .B1(new_n1208), .B2(new_n1174), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT63), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1197), .B1(new_n1174), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT126), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1172), .B(new_n1170), .C1(new_n1206), .C2(new_n1157), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1188), .B2(KEYINPUT63), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT126), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(new_n1211), .A3(new_n1216), .A4(KEYINPUT61), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1203), .B1(new_n1213), .B2(new_n1217), .ZN(G405));
  OAI21_X1  g1018(.A(new_n1206), .B1(new_n1060), .B2(new_n1186), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(new_n1171), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(new_n1198), .ZN(G402));
endmodule


