//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(G146), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  INV_X1    g016(.A(new_n198), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n200), .B1(new_n205), .B2(new_n199), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G110), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT24), .B(G110), .Z(new_n208));
  OR3_X1    g022(.A1(new_n198), .A2(new_n202), .A3(KEYINPUT71), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT71), .B1(new_n198), .B2(new_n202), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI221_X1 g025(.A(new_n193), .B1(G146), .B2(new_n196), .C1(new_n207), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(G110), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n210), .A3(new_n208), .ZN(new_n214));
  INV_X1    g028(.A(new_n193), .ZN(new_n215));
  AOI21_X1  g029(.A(G146), .B1(new_n189), .B2(new_n192), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n219), .B(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n212), .B2(new_n217), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n187), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(G234), .B2(new_n187), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n230), .B(new_n187), .C1(new_n223), .C2(new_n225), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n223), .A2(new_n225), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n229), .A2(G902), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT73), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G472), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G143), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  OR3_X1    g065(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(G146), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n251), .B1(new_n256), .B2(new_n246), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G134), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(KEYINPUT65), .A3(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n260), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT66), .A3(G131), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G131), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n266), .A2(G131), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n257), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n274));
  OAI211_X1 g088(.A(G128), .B(new_n274), .C1(new_n248), .C2(new_n250), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n254), .B(new_n255), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n259), .A2(G134), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n262), .A2(G137), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n277), .B(new_n280), .C1(G131), .C2(new_n266), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n272), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n273), .B1(new_n272), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n245), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G101), .ZN(new_n285));
  NOR2_X1   g099(.A1(G237), .A2(G953), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G210), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n285), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g104(.A(new_n245), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n272), .A2(new_n291), .A3(new_n281), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n272), .A2(new_n294), .A3(new_n291), .A4(new_n281), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n284), .A2(new_n290), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT69), .B1(new_n296), .B2(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(KEYINPUT31), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n293), .A2(new_n295), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n290), .A4(new_n284), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n272), .A2(new_n281), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n245), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n293), .A2(new_n295), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n308), .B2(KEYINPUT28), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n302), .A2(KEYINPUT69), .B1(new_n309), .B2(new_n290), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n238), .B(new_n187), .C1(new_n299), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT32), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n304), .ZN(new_n314));
  INV_X1    g128(.A(new_n290), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n306), .A2(KEYINPUT30), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n272), .A2(new_n273), .A3(new_n281), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n291), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n293), .A2(new_n295), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n301), .A4(new_n290), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n316), .A2(new_n297), .A3(new_n323), .A4(new_n298), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT32), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n238), .A4(new_n187), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n312), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT70), .A2(KEYINPUT29), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n309), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n290), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n315), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n332), .B(new_n187), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G472), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n237), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT99), .ZN(new_n337));
  INV_X1    g151(.A(G116), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G122), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n338), .A2(G122), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n341), .B2(KEYINPUT14), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(KEYINPUT14), .B2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G107), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G128), .B(G143), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(new_n262), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT97), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT13), .B1(new_n247), .B2(G128), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n247), .A2(G128), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT94), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT13), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT95), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n201), .A2(G143), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT13), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT94), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  OAI21_X1  g174(.A(G134), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT96), .B(G134), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n340), .A2(new_n339), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G107), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n346), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n347), .A2(new_n262), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n350), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT97), .B(new_n370), .C1(new_n363), .C2(new_n364), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n349), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n375), .A2(new_n228), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n364), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n354), .B1(new_n201), .B2(G143), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(new_n356), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n382), .A2(new_n353), .A3(new_n355), .A4(new_n358), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT96), .B1(new_n383), .B2(G134), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n371), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT97), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n365), .A2(new_n350), .A3(new_n371), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n349), .A3(new_n376), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT98), .B1(new_n390), .B2(new_n187), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT98), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n392), .B(G902), .C1(new_n378), .C2(new_n389), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G478), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT15), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n337), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n376), .B1(new_n388), .B2(new_n349), .ZN(new_n398));
  INV_X1    g212(.A(new_n349), .ZN(new_n399));
  AOI211_X1 g213(.A(new_n377), .B(new_n399), .C1(new_n386), .C2(new_n387), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n187), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n392), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT98), .B(new_n187), .C1(new_n398), .C2(new_n400), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(new_n337), .A3(new_n396), .A4(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n401), .A2(new_n396), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT100), .B1(new_n397), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n396), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT99), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT100), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n404), .A4(new_n405), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n188), .A2(new_n414), .A3(KEYINPUT19), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(new_n188), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n249), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n286), .A2(G143), .A3(G214), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G143), .B1(new_n286), .B2(G214), .ZN(new_n421));
  OAI21_X1  g235(.A(G131), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n421), .ZN(new_n423));
  INV_X1    g237(.A(G131), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n419), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT90), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n426), .A3(new_n193), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT90), .B1(new_n422), .B2(new_n425), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n188), .B2(new_n249), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n196), .A2(KEYINPUT88), .A3(G146), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT88), .B1(new_n196), .B2(G146), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT87), .B1(new_n196), .B2(G146), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n188), .B2(new_n249), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n438), .A3(new_n432), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT18), .A2(G131), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n423), .A2(new_n419), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n423), .B2(new_n419), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT89), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n440), .A2(new_n447), .A3(new_n444), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n429), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  INV_X1    g264(.A(G104), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n413), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n448), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n447), .B1(new_n440), .B2(new_n444), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n454), .A2(new_n455), .B1(new_n428), .B2(new_n427), .ZN(new_n456));
  INV_X1    g270(.A(new_n452), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT92), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n446), .A2(new_n448), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n215), .A2(new_n216), .ZN(new_n460));
  OAI211_X1 g274(.A(KEYINPUT17), .B(G131), .C1(new_n420), .C2(new_n421), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n422), .A2(new_n425), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n460), .B(new_n461), .C1(KEYINPUT17), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n452), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT20), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n459), .A2(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(KEYINPUT93), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G902), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n468), .A2(new_n470), .B1(G475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(G234), .A2(G237), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n478), .A2(G952), .A3(new_n220), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n478), .A2(G902), .A3(G953), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(G898), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G214), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT3), .B1(new_n451), .B2(G107), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n345), .A3(G104), .ZN(new_n492));
  INV_X1    g306(.A(G101), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n451), .A2(G107), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n345), .A2(G104), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n451), .A2(G107), .ZN(new_n497));
  OAI21_X1  g311(.A(G101), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n197), .A3(G116), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT80), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n501), .A2(new_n197), .A3(KEYINPUT80), .A4(G116), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(G113), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n506), .A3(new_n244), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT81), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT81), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n499), .A2(new_n506), .A3(new_n509), .A4(new_n244), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT79), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G101), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n245), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(G101), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n512), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(new_n245), .A3(new_n512), .A4(new_n515), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n511), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G110), .B(G122), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n523), .B(new_n511), .C1(new_n519), .C2(new_n521), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(KEYINPUT6), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G224), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(G953), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n275), .A2(new_n276), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT82), .A3(new_n194), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT82), .B1(new_n530), .B2(new_n194), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n257), .A2(new_n194), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  INV_X1    g351(.A(new_n529), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n532), .C2(new_n533), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT6), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n522), .A2(new_n541), .A3(new_n524), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n527), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n539), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n523), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n506), .A2(new_n244), .ZN(new_n547));
  INV_X1    g361(.A(new_n499), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT83), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n507), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT83), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT84), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT84), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT85), .B1(new_n532), .B2(new_n533), .ZN(new_n557));
  INV_X1    g371(.A(new_n533), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT85), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n531), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n535), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT86), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n529), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n526), .B(new_n556), .C1(new_n561), .C2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n187), .B1(new_n554), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n489), .B1(new_n543), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n566), .ZN(new_n569));
  AOI22_X1  g383(.A1(KEYINPUT7), .A2(new_n544), .B1(new_n552), .B2(KEYINPUT84), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n527), .A2(new_n540), .A3(new_n542), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n187), .A4(new_n488), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n487), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G469), .ZN(new_n575));
  XOR2_X1   g389(.A(G110), .B(G140), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT75), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n220), .A2(G227), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n277), .A2(new_n499), .A3(KEYINPUT76), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n275), .A2(new_n495), .A3(new_n498), .A4(new_n276), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n518), .A2(new_n257), .A3(new_n515), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n277), .A2(new_n499), .A3(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n581), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT78), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n581), .C1(new_n587), .C2(new_n590), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n596), .A2(new_n580), .A3(new_n589), .A4(new_n588), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n579), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n582), .B(new_n586), .C1(new_n277), .C2(new_n499), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n599), .A2(new_n581), .A3(KEYINPUT12), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT12), .B1(new_n599), .B2(new_n581), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n579), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n575), .B(new_n187), .C1(new_n598), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(G469), .A2(G902), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n597), .A2(KEYINPUT77), .A3(new_n579), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n595), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n611));
  INV_X1    g425(.A(new_n579), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n605), .B(new_n606), .C1(new_n575), .C2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT74), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n574), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n336), .A2(new_n412), .A3(new_n485), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  INV_X1    g436(.A(new_n311), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n238), .B1(new_n324), .B2(new_n187), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n615), .A2(new_n618), .ZN(new_n626));
  INV_X1    g440(.A(new_n237), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n630), .B(new_n633), .C1(new_n398), .C2(new_n400), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n378), .A2(new_n631), .A3(new_n389), .A4(new_n632), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(G478), .A3(new_n187), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n402), .A2(new_n395), .A3(new_n403), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n476), .A2(G475), .ZN(new_n640));
  INV_X1    g454(.A(new_n470), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n573), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n569), .B2(new_n570), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n488), .B1(new_n646), .B2(new_n572), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n483), .B(new_n486), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n629), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT34), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G104), .ZN(G6));
  AOI211_X1 g467(.A(new_n482), .B(new_n487), .C1(new_n568), .C2(new_n573), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n407), .A2(new_n411), .A3(new_n477), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n629), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  NOR2_X1   g472(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n218), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n235), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n232), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n623), .A2(new_n624), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n412), .A2(new_n485), .A3(new_n620), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n327), .A2(new_n335), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n574), .A2(new_n662), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n626), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n479), .B1(new_n480), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n407), .A2(new_n411), .A3(new_n477), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n201), .ZN(G30));
  XOR2_X1   g491(.A(new_n673), .B(KEYINPUT39), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n626), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT40), .Z(new_n680));
  AND3_X1   g494(.A1(new_n407), .A2(new_n411), .A3(new_n643), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n308), .A2(new_n315), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n296), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n327), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n645), .A2(new_n647), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT38), .B1(new_n645), .B2(new_n647), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n487), .B(new_n662), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n680), .A2(new_n681), .A3(new_n685), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  AND3_X1   g506(.A1(new_n639), .A2(new_n643), .A3(new_n674), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n668), .A2(new_n626), .A3(new_n670), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  AOI22_X1  g509(.A1(new_n312), .A2(new_n326), .B1(new_n334), .B2(G472), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n187), .B1(new_n598), .B2(new_n604), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G469), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n618), .A3(new_n605), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n237), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n649), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n655), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NOR2_X1   g519(.A1(new_n696), .A2(new_n669), .ZN(new_n706));
  INV_X1    g520(.A(new_n699), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n412), .A3(new_n485), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n624), .B1(new_n623), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n311), .A2(KEYINPUT103), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n712), .A3(new_n627), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n324), .A2(new_n187), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G472), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n324), .A2(new_n710), .A3(new_n238), .A4(new_n187), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n716), .A3(new_n627), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n648), .A2(new_n699), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n407), .A2(new_n721), .A3(new_n411), .A4(new_n643), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  AND3_X1   g538(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n686), .A2(new_n699), .A3(new_n487), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n693), .A4(new_n662), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  AND3_X1   g542(.A1(new_n568), .A2(new_n486), .A3(new_n573), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n613), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n611), .A2(KEYINPUT105), .A3(new_n612), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n610), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n605), .A2(new_n734), .A3(new_n606), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n730), .A3(new_n618), .A4(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n568), .A2(new_n618), .A3(new_n486), .A4(new_n573), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n605), .A2(new_n734), .A3(new_n606), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT106), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n336), .A2(new_n740), .A3(new_n693), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n336), .A2(new_n740), .A3(KEYINPUT42), .A4(new_n693), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND2_X1  g560(.A1(new_n336), .A2(new_n740), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n675), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n262), .ZN(G36));
  NAND2_X1  g563(.A1(new_n639), .A2(new_n477), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n625), .A2(new_n663), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT44), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n729), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n614), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n732), .A2(KEYINPUT45), .A3(new_n610), .A4(new_n733), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n758), .A3(G469), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n606), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n605), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT46), .B1(new_n759), .B2(new_n606), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n618), .A3(new_n678), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT107), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(new_n766), .A3(new_n618), .A4(new_n678), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n752), .A2(new_n753), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n755), .A2(new_n765), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NAND2_X1  g586(.A1(new_n763), .A2(new_n618), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n618), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n237), .A2(new_n696), .A3(new_n693), .A4(new_n729), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n752), .A2(new_n479), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n698), .A2(new_n605), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n737), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n752), .A2(new_n479), .A3(new_n784), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n781), .B1(new_n789), .B2(new_n336), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n336), .ZN(new_n792));
  AOI211_X1 g606(.A(KEYINPUT116), .B(new_n792), .C1(new_n785), .C2(new_n788), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n794), .A3(KEYINPUT48), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n688), .A2(new_n689), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n486), .A3(new_n699), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n782), .A2(new_n720), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n685), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n627), .A3(new_n479), .A4(new_n784), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n643), .A3(new_n639), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n716), .A2(new_n713), .A3(new_n662), .A4(new_n717), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n789), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n782), .A2(new_n720), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n783), .B(KEYINPUT108), .Z(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n618), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n806), .B(new_n729), .C1(new_n777), .C2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n800), .A2(new_n805), .A3(KEYINPUT51), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT48), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n790), .B2(new_n793), .ZN(new_n812));
  OAI211_X1 g626(.A(G952), .B(new_n220), .C1(new_n802), .C2(new_n644), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n806), .B2(new_n726), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n795), .A2(new_n810), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n800), .A2(new_n805), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n808), .B1(new_n777), .B2(KEYINPUT114), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(KEYINPUT114), .B2(new_n777), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n729), .A3(new_n806), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n694), .B(new_n727), .C1(new_n671), .C2(new_n675), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT110), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n617), .A2(new_n673), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n735), .A2(new_n663), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n232), .A2(new_n661), .A3(new_n825), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT110), .B1(new_n738), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n826), .A2(new_n828), .B1(new_n327), .B2(new_n684), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n681), .A2(new_n829), .A3(new_n830), .A4(new_n574), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n826), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n685), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n407), .A2(new_n411), .A3(new_n643), .A4(new_n574), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT111), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n823), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n823), .A2(new_n836), .A3(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n644), .B2(new_n648), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n468), .A2(new_n470), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n844), .A2(new_n640), .B1(new_n637), .B2(new_n638), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(KEYINPUT109), .A3(new_n654), .ZN(new_n846));
  INV_X1    g660(.A(new_n406), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n643), .B1(new_n847), .B2(new_n409), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n843), .A2(new_n846), .B1(new_n848), .B2(new_n654), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n621), .B(new_n665), .C1(new_n849), .C2(new_n628), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n409), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n662), .A2(new_n674), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n568), .A2(new_n486), .A3(new_n573), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n853), .A2(new_n643), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n852), .A2(new_n668), .A3(new_n626), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n740), .A2(new_n804), .A3(new_n693), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n856), .B(new_n857), .C1(new_n747), .C2(new_n675), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n700), .B1(new_n655), .B2(new_n649), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n745), .A2(new_n708), .A3(new_n723), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n841), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n745), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n723), .A3(new_n708), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n850), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n823), .A2(new_n836), .A3(KEYINPUT52), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(new_n823), .B2(new_n836), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n866), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n869), .A2(new_n870), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n850), .A2(new_n858), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n867), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT112), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n865), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n864), .B1(new_n878), .B2(new_n865), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n841), .A2(new_n868), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n873), .A2(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n821), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n807), .B(KEYINPUT49), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n627), .A2(new_n618), .A3(new_n486), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n796), .A2(new_n750), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n801), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(G75));
  NAND2_X1  g704(.A1(new_n877), .A2(new_n881), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(G210), .A3(G902), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n527), .A2(new_n542), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT117), .Z(new_n895));
  XNOR2_X1  g709(.A(new_n540), .B(KEYINPUT55), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n892), .A2(new_n893), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n892), .B2(new_n893), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n220), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  XOR2_X1   g716(.A(new_n606), .B(KEYINPUT57), .Z(new_n903));
  AND3_X1   g717(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n882), .B1(new_n877), .B2(new_n881), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n598), .B2(new_n604), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n891), .A2(G902), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(new_n759), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n901), .B1(new_n907), .B2(new_n909), .ZN(G54));
  INV_X1    g724(.A(new_n465), .ZN(new_n911));
  NAND2_X1  g725(.A1(KEYINPUT58), .A2(G475), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n901), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(G60));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n873), .B2(new_n883), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n920), .B2(new_n636), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n634), .B2(new_n635), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n904), .B2(new_n905), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT119), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n925), .B(new_n922), .C1(new_n904), .C2(new_n905), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n877), .B2(new_n881), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n930), .A2(KEYINPUT120), .A3(new_n233), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT120), .B1(new_n930), .B2(new_n233), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n930), .B2(new_n660), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n930), .A2(new_n660), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n914), .B1(new_n930), .B2(new_n233), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(G66));
  NOR3_X1   g754(.A1(new_n481), .A2(new_n528), .A3(new_n220), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n865), .A2(new_n850), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n220), .ZN(new_n943));
  INV_X1    g757(.A(new_n895), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(G898), .B2(new_n220), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n792), .A2(new_n679), .A3(new_n854), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT123), .B(new_n644), .C1(new_n852), .C2(new_n643), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n848), .B2(new_n845), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n771), .A2(new_n779), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n691), .B1(KEYINPUT122), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT121), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n822), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n953), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n955), .B2(new_n957), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n220), .ZN(new_n963));
  NAND3_X1  g777(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n282), .A2(new_n283), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(new_n417), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n748), .B1(new_n777), .B2(new_n778), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n792), .A2(new_n834), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n765), .A2(new_n767), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n771), .A2(new_n970), .A3(new_n745), .A4(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n220), .B1(new_n973), .B2(new_n957), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n672), .A2(new_n220), .A3(G227), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n968), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n947), .B1(new_n969), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(KEYINPUT124), .B(new_n977), .C1(new_n965), .C2(new_n968), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G72));
  OAI21_X1  g795(.A(new_n290), .B1(new_n319), .B2(new_n320), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n961), .A2(new_n942), .A3(new_n962), .ZN(new_n983));
  XNOR2_X1  g797(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n987), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n973), .A2(new_n957), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n942), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n914), .B1(new_n991), .B2(new_n333), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n333), .A2(new_n982), .A3(new_n986), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT127), .Z(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n877), .B2(new_n871), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n988), .A2(new_n992), .A3(new_n995), .ZN(G57));
endmodule


