

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G168), .A2(n599), .ZN(n600) );
  XNOR2_X1 U550 ( .A(n613), .B(KEYINPUT13), .ZN(n614) );
  XNOR2_X1 U551 ( .A(n543), .B(KEYINPUT64), .ZN(n874) );
  NOR2_X1 U552 ( .A1(n663), .A2(n596), .ZN(n514) );
  NOR2_X1 U553 ( .A1(n689), .A2(n675), .ZN(n515) );
  INV_X1 U554 ( .A(G8), .ZN(n596) );
  AND2_X1 U555 ( .A1(n664), .A2(n514), .ZN(n598) );
  INV_X1 U556 ( .A(KEYINPUT90), .ZN(n594) );
  AND2_X1 U557 ( .A1(n749), .A2(G40), .ZN(n714) );
  INV_X1 U558 ( .A(G2105), .ZN(n542) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XNOR2_X1 U560 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X1 U561 ( .A1(G651), .A2(n524), .ZN(n776) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n779) );
  NAND2_X1 U563 ( .A1(n779), .A2(G89), .ZN(n516) );
  XNOR2_X1 U564 ( .A(n516), .B(KEYINPUT4), .ZN(n520) );
  XNOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .ZN(n517) );
  XNOR2_X1 U566 ( .A(n517), .B(KEYINPUT67), .ZN(n524) );
  INV_X1 U567 ( .A(G651), .ZN(n522) );
  OR2_X1 U568 ( .A1(n524), .A2(n522), .ZN(n518) );
  XOR2_X2 U569 ( .A(KEYINPUT68), .B(n518), .Z(n780) );
  NAND2_X1 U570 ( .A1(G76), .A2(n780), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n521), .B(KEYINPUT5), .ZN(n529) );
  NOR2_X1 U573 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n523), .Z(n775) );
  NAND2_X1 U575 ( .A1(G63), .A2(n775), .ZN(n526) );
  NAND2_X1 U576 ( .A1(G51), .A2(n776), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U578 ( .A(KEYINPUT6), .B(n527), .Z(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U581 ( .A1(G48), .A2(n776), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G86), .A2(n779), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n780), .A2(G73), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT2), .B(n533), .Z(n534) );
  NOR2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n775), .A2(G61), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(G305) );
  XOR2_X2 U589 ( .A(KEYINPUT17), .B(n538), .Z(n869) );
  NAND2_X1 U590 ( .A1(G138), .A2(n869), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n542), .A2(G2104), .ZN(n539) );
  XNOR2_X2 U592 ( .A(n539), .B(KEYINPUT65), .ZN(n870) );
  NAND2_X1 U593 ( .A1(G102), .A2(n870), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n547) );
  AND2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U596 ( .A1(n873), .A2(G114), .ZN(n545) );
  NOR2_X1 U597 ( .A1(n542), .A2(G2104), .ZN(n543) );
  NAND2_X1 U598 ( .A1(G126), .A2(n874), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U600 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U601 ( .A1(G49), .A2(n776), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G87), .A2(n524), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n775), .A2(n550), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G651), .A2(G74), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(G288) );
  NAND2_X1 U607 ( .A1(n776), .A2(G52), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n775), .A2(G64), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U610 ( .A1(G90), .A2(n779), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G77), .A2(n780), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U613 ( .A(n557), .B(KEYINPUT9), .ZN(n558) );
  XNOR2_X1 U614 ( .A(n558), .B(KEYINPUT71), .ZN(n559) );
  NOR2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U616 ( .A(KEYINPUT72), .B(n561), .Z(G301) );
  INV_X1 U617 ( .A(G301), .ZN(G171) );
  NAND2_X1 U618 ( .A1(n779), .A2(G91), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G78), .A2(n780), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U621 ( .A(KEYINPUT73), .B(n564), .ZN(n568) );
  NAND2_X1 U622 ( .A1(G65), .A2(n775), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G53), .A2(n776), .ZN(n565) );
  AND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(G299) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G62), .A2(n775), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G88), .A2(n779), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G75), .A2(n780), .ZN(n571) );
  XNOR2_X1 U631 ( .A(KEYINPUT79), .B(n571), .ZN(n572) );
  NOR2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n776), .A2(G50), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n575), .A2(n574), .ZN(G303) );
  NAND2_X1 U635 ( .A1(G72), .A2(n780), .ZN(n576) );
  XOR2_X1 U636 ( .A(KEYINPUT69), .B(n576), .Z(n578) );
  NAND2_X1 U637 ( .A1(n779), .A2(G85), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U639 ( .A(KEYINPUT70), .B(n579), .Z(n583) );
  NAND2_X1 U640 ( .A1(G60), .A2(n775), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G47), .A2(n776), .ZN(n580) );
  AND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(G290) );
  XOR2_X1 U644 ( .A(G1981), .B(G305), .Z(n948) );
  NAND2_X1 U645 ( .A1(G101), .A2(n870), .ZN(n584) );
  XNOR2_X1 U646 ( .A(KEYINPUT23), .B(n584), .ZN(n591) );
  NAND2_X1 U647 ( .A1(G137), .A2(n869), .ZN(n585) );
  XNOR2_X1 U648 ( .A(n585), .B(KEYINPUT66), .ZN(n589) );
  NAND2_X1 U649 ( .A1(G125), .A2(n874), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n873), .A2(G113), .ZN(n586) );
  AND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U653 ( .A1(n591), .A2(n590), .ZN(n749) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NAND2_X2 U655 ( .A1(n714), .A2(n715), .ZN(n655) );
  NAND2_X1 U656 ( .A1(G8), .A2(n655), .ZN(n689) );
  NOR2_X1 U657 ( .A1(G1976), .A2(G288), .ZN(n673) );
  INV_X1 U658 ( .A(n673), .ZN(n938) );
  NOR2_X1 U659 ( .A1(n689), .A2(n938), .ZN(n592) );
  NAND2_X1 U660 ( .A1(KEYINPUT33), .A2(n592), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n948), .A2(n593), .ZN(n679) );
  NOR2_X1 U662 ( .A1(G1966), .A2(n689), .ZN(n595) );
  XNOR2_X1 U663 ( .A(n595), .B(n594), .ZN(n664) );
  NOR2_X1 U664 ( .A1(G2084), .A2(n655), .ZN(n663) );
  XOR2_X1 U665 ( .A(KEYINPUT92), .B(KEYINPUT30), .Z(n597) );
  XNOR2_X1 U666 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT93), .ZN(n604) );
  INV_X1 U668 ( .A(G1961), .ZN(n925) );
  NAND2_X1 U669 ( .A1(n655), .A2(n925), .ZN(n602) );
  INV_X1 U670 ( .A(n655), .ZN(n639) );
  XNOR2_X1 U671 ( .A(G2078), .B(KEYINPUT25), .ZN(n962) );
  NAND2_X1 U672 ( .A1(n639), .A2(n962), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n607) );
  OR2_X1 U674 ( .A1(n607), .A2(G171), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT31), .B(KEYINPUT94), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n653) );
  NAND2_X1 U678 ( .A1(n607), .A2(G171), .ZN(n651) );
  NAND2_X1 U679 ( .A1(n775), .A2(G56), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT14), .B(n608), .Z(n617) );
  NAND2_X1 U681 ( .A1(n779), .A2(G81), .ZN(n609) );
  XNOR2_X1 U682 ( .A(KEYINPUT12), .B(n609), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G68), .A2(n780), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT76), .ZN(n611) );
  AND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n615) );
  INV_X1 U686 ( .A(KEYINPUT77), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n776), .A2(G43), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n932) );
  INV_X1 U690 ( .A(G1996), .ZN(n965) );
  NOR2_X1 U691 ( .A1(n655), .A2(n965), .ZN(n620) );
  XOR2_X1 U692 ( .A(n620), .B(KEYINPUT26), .Z(n622) );
  NAND2_X1 U693 ( .A1(n655), .A2(G1341), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U695 ( .A1(n932), .A2(n623), .ZN(n636) );
  NAND2_X1 U696 ( .A1(G66), .A2(n775), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G79), .A2(n780), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G54), .A2(n776), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G92), .A2(n779), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U703 ( .A(KEYINPUT15), .B(n630), .Z(n884) );
  NAND2_X1 U704 ( .A1(n636), .A2(n884), .ZN(n635) );
  INV_X1 U705 ( .A(G2067), .ZN(n963) );
  NOR2_X1 U706 ( .A1(n655), .A2(n963), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT91), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n655), .A2(G1348), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n638) );
  OR2_X1 U711 ( .A1(n884), .A2(n636), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n644) );
  INV_X1 U713 ( .A(G299), .ZN(n935) );
  NAND2_X1 U714 ( .A1(n639), .A2(G2072), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(KEYINPUT27), .ZN(n642) );
  AND2_X1 U716 ( .A1(G1956), .A2(n655), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n935), .A2(n645), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n935), .A2(n645), .ZN(n646) );
  XOR2_X1 U721 ( .A(n646), .B(KEYINPUT28), .Z(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U723 ( .A(KEYINPUT29), .B(n649), .Z(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n665) );
  NAND2_X1 U726 ( .A1(n665), .A2(G286), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n654), .B(KEYINPUT96), .ZN(n660) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n689), .ZN(n657) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n655), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n658), .A2(G303), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n661), .A2(G8), .ZN(n662) );
  XNOR2_X1 U734 ( .A(KEYINPUT32), .B(n662), .ZN(n670) );
  NAND2_X1 U735 ( .A1(G8), .A2(n663), .ZN(n668) );
  AND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT95), .B(n666), .Z(n667) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n687) );
  NOR2_X1 U740 ( .A1(G1971), .A2(G303), .ZN(n671) );
  XOR2_X1 U741 ( .A(n671), .B(KEYINPUT97), .Z(n672) );
  NOR2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n687), .A2(n674), .ZN(n676) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n937) );
  INV_X1 U745 ( .A(n937), .ZN(n675) );
  AND2_X1 U746 ( .A1(n676), .A2(n515), .ZN(n677) );
  NOR2_X1 U747 ( .A1(KEYINPUT33), .A2(n677), .ZN(n678) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n684) );
  NOR2_X1 U749 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(KEYINPUT89), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n681), .B(KEYINPUT24), .ZN(n682) );
  NOR2_X1 U752 ( .A1(n682), .A2(n689), .ZN(n683) );
  NOR2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n721) );
  NOR2_X1 U754 ( .A1(G2090), .A2(G303), .ZN(n685) );
  NAND2_X1 U755 ( .A1(G8), .A2(n685), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n686), .B(KEYINPUT98), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n719) );
  NAND2_X1 U759 ( .A1(G117), .A2(n873), .ZN(n692) );
  NAND2_X1 U760 ( .A1(G141), .A2(n869), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n698) );
  NAND2_X1 U762 ( .A1(G105), .A2(n870), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT88), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(KEYINPUT38), .ZN(n696) );
  NAND2_X1 U765 ( .A1(G129), .A2(n874), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n855) );
  AND2_X1 U768 ( .A1(n965), .A2(n855), .ZN(n699) );
  XOR2_X1 U769 ( .A(KEYINPUT99), .B(n699), .Z(n983) );
  NAND2_X1 U770 ( .A1(G107), .A2(n873), .ZN(n701) );
  NAND2_X1 U771 ( .A1(G131), .A2(n869), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G95), .A2(n870), .ZN(n702) );
  XOR2_X1 U774 ( .A(KEYINPUT87), .B(n702), .Z(n704) );
  NAND2_X1 U775 ( .A1(G119), .A2(n874), .ZN(n703) );
  NAND2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n846) );
  INV_X1 U778 ( .A(G1991), .ZN(n959) );
  NOR2_X1 U779 ( .A1(n846), .A2(n959), .ZN(n708) );
  NOR2_X1 U780 ( .A1(n855), .A2(n965), .ZN(n707) );
  NOR2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n723) );
  INV_X1 U782 ( .A(n723), .ZN(n992) );
  NOR2_X1 U783 ( .A1(G1986), .A2(G290), .ZN(n709) );
  AND2_X1 U784 ( .A1(n959), .A2(n846), .ZN(n991) );
  NOR2_X1 U785 ( .A1(n709), .A2(n991), .ZN(n710) );
  XNOR2_X1 U786 ( .A(n710), .B(KEYINPUT100), .ZN(n711) );
  NOR2_X1 U787 ( .A1(n992), .A2(n711), .ZN(n712) );
  NOR2_X1 U788 ( .A1(n983), .A2(n712), .ZN(n713) );
  XNOR2_X1 U789 ( .A(KEYINPUT39), .B(n713), .ZN(n718) );
  INV_X1 U790 ( .A(n714), .ZN(n716) );
  NOR2_X1 U791 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U792 ( .A(n717), .B(KEYINPUT84), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n718), .A2(n744), .ZN(n722) );
  AND2_X1 U794 ( .A1(n719), .A2(n722), .ZN(n720) );
  NAND2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n728) );
  INV_X1 U796 ( .A(n722), .ZN(n726) );
  XOR2_X1 U797 ( .A(G1986), .B(G290), .Z(n952) );
  NAND2_X1 U798 ( .A1(n952), .A2(n723), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n724), .A2(n744), .ZN(n725) );
  OR2_X1 U800 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n741) );
  NAND2_X1 U802 ( .A1(G140), .A2(n869), .ZN(n730) );
  NAND2_X1 U803 ( .A1(G104), .A2(n870), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n732) );
  XOR2_X1 U805 ( .A(KEYINPUT85), .B(KEYINPUT34), .Z(n731) );
  XNOR2_X1 U806 ( .A(n732), .B(n731), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n873), .A2(G116), .ZN(n734) );
  NAND2_X1 U808 ( .A1(G128), .A2(n874), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n736) );
  XOR2_X1 U810 ( .A(KEYINPUT35), .B(KEYINPUT86), .Z(n735) );
  XNOR2_X1 U811 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U813 ( .A(KEYINPUT36), .B(n739), .ZN(n856) );
  XNOR2_X1 U814 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n856), .A2(n742), .ZN(n993) );
  NAND2_X1 U816 ( .A1(n993), .A2(n744), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n741), .A2(n740), .ZN(n746) );
  AND2_X1 U818 ( .A1(n856), .A2(n742), .ZN(n743) );
  XOR2_X1 U819 ( .A(KEYINPUT101), .B(n743), .Z(n1002) );
  NAND2_X1 U820 ( .A1(n1002), .A2(n744), .ZN(n745) );
  NAND2_X1 U821 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U822 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n747) );
  XNOR2_X1 U823 ( .A(n748), .B(n747), .ZN(G329) );
  BUF_X1 U824 ( .A(n749), .Z(G160) );
  AND2_X1 U825 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U826 ( .A(G132), .ZN(G219) );
  INV_X1 U827 ( .A(G82), .ZN(G220) );
  NAND2_X1 U828 ( .A1(G7), .A2(G661), .ZN(n750) );
  XNOR2_X1 U829 ( .A(n750), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U830 ( .A(G223), .ZN(n813) );
  NAND2_X1 U831 ( .A1(n813), .A2(G567), .ZN(n751) );
  XNOR2_X1 U832 ( .A(n751), .B(KEYINPUT11), .ZN(n752) );
  XNOR2_X1 U833 ( .A(KEYINPUT75), .B(n752), .ZN(G234) );
  INV_X1 U834 ( .A(G860), .ZN(n758) );
  OR2_X1 U835 ( .A1(n932), .A2(n758), .ZN(G153) );
  NAND2_X1 U836 ( .A1(G301), .A2(G868), .ZN(n754) );
  INV_X1 U837 ( .A(n884), .ZN(n943) );
  INV_X1 U838 ( .A(G868), .ZN(n755) );
  NAND2_X1 U839 ( .A1(n943), .A2(n755), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(G284) );
  NOR2_X1 U841 ( .A1(G286), .A2(n755), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G868), .A2(G299), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n757), .A2(n756), .ZN(G297) );
  NAND2_X1 U844 ( .A1(n758), .A2(G559), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n759), .A2(n884), .ZN(n760) );
  XNOR2_X1 U846 ( .A(n760), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U847 ( .A1(n884), .A2(G868), .ZN(n761) );
  NOR2_X1 U848 ( .A1(G559), .A2(n761), .ZN(n762) );
  XNOR2_X1 U849 ( .A(n762), .B(KEYINPUT78), .ZN(n764) );
  NOR2_X1 U850 ( .A1(n932), .A2(G868), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(G282) );
  NAND2_X1 U852 ( .A1(G123), .A2(n874), .ZN(n765) );
  XNOR2_X1 U853 ( .A(n765), .B(KEYINPUT18), .ZN(n767) );
  NAND2_X1 U854 ( .A1(G111), .A2(n873), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G135), .A2(n869), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G99), .A2(n870), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n990) );
  XNOR2_X1 U860 ( .A(n990), .B(G2096), .ZN(n773) );
  INV_X1 U861 ( .A(G2100), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(G156) );
  NAND2_X1 U863 ( .A1(n884), .A2(G559), .ZN(n793) );
  XNOR2_X1 U864 ( .A(n932), .B(n793), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n774), .A2(G860), .ZN(n785) );
  NAND2_X1 U866 ( .A1(G67), .A2(n775), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G55), .A2(n776), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n779), .A2(G93), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G80), .A2(n780), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n796) );
  XNOR2_X1 U873 ( .A(n785), .B(n796), .ZN(G145) );
  INV_X1 U874 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U875 ( .A(G166), .B(G305), .ZN(n786) );
  XNOR2_X1 U876 ( .A(n786), .B(G290), .ZN(n789) );
  XOR2_X1 U877 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n787) );
  XNOR2_X1 U878 ( .A(G288), .B(n787), .ZN(n788) );
  XOR2_X1 U879 ( .A(n789), .B(n788), .Z(n791) );
  XNOR2_X1 U880 ( .A(n935), .B(n796), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(n932), .ZN(n885) );
  XNOR2_X1 U883 ( .A(n885), .B(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n794), .A2(G868), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n795), .B(KEYINPUT81), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n796), .A2(G868), .ZN(n797) );
  NOR2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U888 ( .A(KEYINPUT82), .B(n799), .Z(G295) );
  NAND2_X1 U889 ( .A1(G2084), .A2(G2078), .ZN(n800) );
  XNOR2_X1 U890 ( .A(n800), .B(KEYINPUT20), .ZN(n801) );
  XNOR2_X1 U891 ( .A(n801), .B(KEYINPUT83), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n802), .A2(G2090), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(n803), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n804), .A2(G2072), .ZN(G158) );
  XOR2_X1 U895 ( .A(KEYINPUT74), .B(G57), .Z(G237) );
  XNOR2_X1 U896 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U897 ( .A1(G108), .A2(G69), .ZN(n805) );
  NOR2_X1 U898 ( .A1(G237), .A2(n805), .ZN(n806) );
  NAND2_X1 U899 ( .A1(G120), .A2(n806), .ZN(n818) );
  NAND2_X1 U900 ( .A1(n818), .A2(G567), .ZN(n811) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n807) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(n807), .Z(n808) );
  NOR2_X1 U903 ( .A1(G218), .A2(n808), .ZN(n809) );
  NAND2_X1 U904 ( .A1(G96), .A2(n809), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G2106), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n820) );
  NAND2_X1 U907 ( .A1(G483), .A2(G661), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n820), .A2(n812), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n815), .A2(G36), .ZN(G176) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U912 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G1), .A2(G3), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n817), .B(KEYINPUT104), .ZN(G188) );
  XNOR2_X1 U916 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  XNOR2_X1 U917 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  NOR2_X1 U921 ( .A1(n819), .A2(n818), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  INV_X1 U923 ( .A(n820), .ZN(G319) );
  XNOR2_X1 U924 ( .A(G1996), .B(KEYINPUT41), .ZN(n830) );
  XOR2_X1 U925 ( .A(G1991), .B(G1976), .Z(n822) );
  XNOR2_X1 U926 ( .A(G1966), .B(G1981), .ZN(n821) );
  XNOR2_X1 U927 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U928 ( .A(G1986), .B(G1971), .Z(n824) );
  XNOR2_X1 U929 ( .A(G1961), .B(G1956), .ZN(n823) );
  XNOR2_X1 U930 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U931 ( .A(n826), .B(n825), .Z(n828) );
  XNOR2_X1 U932 ( .A(KEYINPUT106), .B(G2474), .ZN(n827) );
  XNOR2_X1 U933 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U934 ( .A(n830), .B(n829), .ZN(G229) );
  XOR2_X1 U935 ( .A(G2100), .B(G2096), .Z(n832) );
  XNOR2_X1 U936 ( .A(KEYINPUT42), .B(G2678), .ZN(n831) );
  XNOR2_X1 U937 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(G2090), .Z(n834) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U940 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U941 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U942 ( .A(G2084), .B(G2078), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n838), .B(n837), .ZN(G227) );
  NAND2_X1 U944 ( .A1(G124), .A2(n874), .ZN(n839) );
  XNOR2_X1 U945 ( .A(n839), .B(KEYINPUT44), .ZN(n841) );
  NAND2_X1 U946 ( .A1(G112), .A2(n873), .ZN(n840) );
  NAND2_X1 U947 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U948 ( .A1(G136), .A2(n869), .ZN(n843) );
  NAND2_X1 U949 ( .A1(G100), .A2(n870), .ZN(n842) );
  NAND2_X1 U950 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U951 ( .A1(n845), .A2(n844), .ZN(G162) );
  XNOR2_X1 U952 ( .A(G164), .B(n846), .ZN(n853) );
  XOR2_X1 U953 ( .A(KEYINPUT110), .B(KEYINPUT108), .Z(n848) );
  XNOR2_X1 U954 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n847) );
  XNOR2_X1 U955 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U956 ( .A(n849), .B(KEYINPUT112), .Z(n851) );
  XNOR2_X1 U957 ( .A(n990), .B(KEYINPUT48), .ZN(n850) );
  XNOR2_X1 U958 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U959 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U960 ( .A(n854), .B(G162), .Z(n858) );
  XOR2_X1 U961 ( .A(n856), .B(n855), .Z(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n868) );
  NAND2_X1 U963 ( .A1(n873), .A2(G118), .ZN(n860) );
  NAND2_X1 U964 ( .A1(G130), .A2(n874), .ZN(n859) );
  NAND2_X1 U965 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n869), .A2(G142), .ZN(n861) );
  XOR2_X1 U967 ( .A(KEYINPUT107), .B(n861), .Z(n863) );
  NAND2_X1 U968 ( .A1(n870), .A2(G106), .ZN(n862) );
  NAND2_X1 U969 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U970 ( .A(n864), .B(KEYINPUT45), .Z(n865) );
  NOR2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U972 ( .A(n868), .B(n867), .Z(n882) );
  NAND2_X1 U973 ( .A1(G139), .A2(n869), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G103), .A2(n870), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U976 ( .A1(n873), .A2(G115), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G127), .A2(n874), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n877), .ZN(n878) );
  XNOR2_X1 U980 ( .A(KEYINPUT109), .B(n878), .ZN(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n985) );
  XNOR2_X1 U982 ( .A(n985), .B(G160), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U984 ( .A1(G37), .A2(n883), .ZN(G395) );
  XNOR2_X1 U985 ( .A(n884), .B(G286), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n887), .B(G301), .ZN(n888) );
  NOR2_X1 U988 ( .A1(G37), .A2(n888), .ZN(G397) );
  XOR2_X1 U989 ( .A(KEYINPUT103), .B(G2427), .Z(n890) );
  XNOR2_X1 U990 ( .A(G2435), .B(G2438), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n897) );
  XOR2_X1 U992 ( .A(G2443), .B(G2430), .Z(n892) );
  XNOR2_X1 U993 ( .A(G2454), .B(G2446), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U995 ( .A(n893), .B(G2451), .Z(n895) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n898), .A2(G14), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n904), .ZN(n901) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n899) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n899), .ZN(n900) );
  NOR2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n903) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(n904), .ZN(G401) );
  XNOR2_X1 U1008 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1015) );
  XOR2_X1 U1009 ( .A(G1986), .B(G24), .Z(n908) );
  XNOR2_X1 U1010 ( .A(G1971), .B(G22), .ZN(n906) );
  XNOR2_X1 U1011 ( .A(G23), .B(G1976), .ZN(n905) );
  NOR2_X1 U1012 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1013 ( .A1(n908), .A2(n907), .ZN(n910) );
  XNOR2_X1 U1014 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n909) );
  XNOR2_X1 U1015 ( .A(n910), .B(n909), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT59), .ZN(n911) );
  XNOR2_X1 U1017 ( .A(n911), .B(G4), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n913) );
  XNOR2_X1 U1019 ( .A(G1981), .B(G6), .ZN(n912) );
  NOR2_X1 U1020 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1021 ( .A1(n915), .A2(n914), .ZN(n918) );
  XOR2_X1 U1022 ( .A(G20), .B(G1956), .Z(n916) );
  XNOR2_X1 U1023 ( .A(KEYINPUT123), .B(n916), .ZN(n917) );
  NOR2_X1 U1024 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1025 ( .A(n919), .B(KEYINPUT60), .Z(n920) );
  XNOR2_X1 U1026 ( .A(KEYINPUT124), .B(n920), .ZN(n922) );
  XNOR2_X1 U1027 ( .A(G21), .B(G1966), .ZN(n921) );
  NOR2_X1 U1028 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1029 ( .A1(n924), .A2(n923), .ZN(n928) );
  XOR2_X1 U1030 ( .A(G5), .B(n925), .Z(n926) );
  XNOR2_X1 U1031 ( .A(KEYINPUT122), .B(n926), .ZN(n927) );
  NOR2_X1 U1032 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1033 ( .A(KEYINPUT61), .B(n929), .Z(n930) );
  NOR2_X1 U1034 ( .A1(G16), .A2(n930), .ZN(n1013) );
  XNOR2_X1 U1035 ( .A(G16), .B(KEYINPUT119), .ZN(n931) );
  XNOR2_X1 U1036 ( .A(n931), .B(KEYINPUT56), .ZN(n957) );
  XNOR2_X1 U1037 ( .A(n932), .B(G1341), .ZN(n934) );
  XNOR2_X1 U1038 ( .A(G301), .B(G1961), .ZN(n933) );
  NOR2_X1 U1039 ( .A1(n934), .A2(n933), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n935), .B(G1956), .ZN(n936) );
  XNOR2_X1 U1041 ( .A(n936), .B(KEYINPUT120), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(G1971), .B(G303), .ZN(n939) );
  NOR2_X1 U1044 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(G1348), .B(n943), .ZN(n944) );
  NOR2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G168), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(n950), .B(KEYINPUT57), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1054 ( .A(KEYINPUT121), .B(n955), .Z(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n1010) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n958) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n958), .ZN(n977) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G35), .ZN(n975) );
  XOR2_X1 U1059 ( .A(G2072), .B(G33), .Z(n961) );
  XNOR2_X1 U1060 ( .A(n959), .B(G25), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G27), .B(n962), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G26), .B(n963), .ZN(n964) );
  NAND2_X1 U1064 ( .A1(n964), .A2(G28), .ZN(n968) );
  XOR2_X1 U1065 ( .A(G32), .B(n965), .Z(n966) );
  XNOR2_X1 U1066 ( .A(KEYINPUT116), .B(n966), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT118), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT117), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(G29), .A2(n980), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT55), .ZN(n1008) );
  XOR2_X1 U1077 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1079 ( .A(KEYINPUT51), .B(n984), .Z(n1004) );
  XOR2_X1 U1080 ( .A(n985), .B(KEYINPUT115), .Z(n986) );
  XOR2_X1 U1081 ( .A(G2072), .B(n986), .Z(n988) );
  XOR2_X1 U1082 ( .A(G164), .B(G2078), .Z(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT50), .B(n989), .ZN(n1000) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1088 ( .A(G2084), .B(G160), .Z(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT114), .B(n996), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT52), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(G29), .A2(n1006), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(G11), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1015), .B(n1014), .ZN(G311) );
  XNOR2_X1 U1101 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

