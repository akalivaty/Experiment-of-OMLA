//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n214), .A2(KEYINPUT65), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(KEYINPUT65), .B2(new_n214), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT67), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT68), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G116), .A2(G270), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n211), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(KEYINPUT69), .ZN(new_n235));
  AND2_X1   g0035(.A1(new_n234), .A2(KEYINPUT69), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n224), .B(new_n237), .C1(new_n235), .C2(new_n233), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT70), .Z(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(KEYINPUT73), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(KEYINPUT10), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n203), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n209), .A2(G33), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n259), .B1(new_n260), .B2(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n215), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(new_n209), .A3(G1), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n208), .B2(G20), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n271), .A2(new_n273), .B1(new_n272), .B2(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n277), .B(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G222), .ZN(new_n284));
  OR2_X1    g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(G1698), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n284), .B1(new_n226), .B2(new_n287), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(new_n292), .A3(G274), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT71), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  INV_X1    g0100(.A(new_n215), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n291), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT71), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n297), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n293), .A2(new_n297), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n299), .A2(new_n304), .B1(new_n305), .B2(G226), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n294), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n294), .B2(new_n306), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n275), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(KEYINPUT9), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n257), .B(new_n258), .C1(new_n279), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n314), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n277), .B(KEYINPUT72), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n256), .A4(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n275), .C1(G179), .C2(new_n307), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n315), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n267), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n209), .A2(G33), .A3(G77), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT76), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n269), .A2(G1), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G20), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n332), .A2(KEYINPUT12), .A3(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT12), .B1(new_n332), .B2(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n325), .B1(new_n208), .B2(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n333), .A2(new_n334), .B1(new_n271), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n329), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT77), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n337), .A2(KEYINPUT77), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n241), .A2(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n287), .B(new_n344), .C1(G226), .C2(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n292), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n299), .A2(new_n304), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n305), .A2(G238), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n348), .A3(new_n350), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n355), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n357), .B(new_n347), .C1(new_n352), .C2(new_n353), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n343), .B(G169), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n355), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(G179), .C1(new_n361), .C2(new_n354), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n353), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n351), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n357), .B1(new_n365), .B2(new_n347), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n360), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n343), .B1(new_n367), .B2(G169), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n342), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n356), .B2(new_n358), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n360), .B(G190), .C1(new_n361), .C2(new_n354), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n338), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n292), .A2(G232), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT80), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n292), .A2(new_n374), .A3(KEYINPUT80), .A4(G232), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n304), .A2(new_n299), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT79), .ZN(new_n381));
  OAI211_X1 g0181(.A(G226), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n382));
  INV_X1    g0182(.A(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(G223), .B(new_n383), .C1(new_n280), .C2(new_n281), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n293), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n379), .A2(G179), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n319), .B1(new_n379), .B2(new_n386), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  INV_X1    g0190(.A(G159), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n262), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  XNOR2_X1  g0194(.A(G58), .B(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(G20), .ZN(new_n396));
  AND2_X1   g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n394), .B(G20), .C1(new_n397), .C2(new_n218), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n393), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n285), .A2(new_n209), .A3(new_n286), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n286), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n325), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n390), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n282), .B2(new_n209), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n280), .A2(new_n281), .A3(new_n402), .A4(G20), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n397), .B2(new_n218), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT78), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n392), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n406), .A2(new_n267), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n264), .B1(new_n208), .B2(G20), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n271), .B1(new_n270), .B2(new_n264), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n389), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(KEYINPUT18), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n389), .B2(new_n417), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n379), .A2(new_n386), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G200), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n379), .A2(G190), .A3(new_n386), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n414), .A2(new_n424), .A3(new_n416), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n283), .A2(G232), .ZN(new_n428));
  INV_X1    g0228(.A(G107), .ZN(new_n429));
  INV_X1    g0229(.A(G238), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n428), .B1(new_n429), .B2(new_n287), .C1(new_n430), .C2(new_n289), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n293), .ZN(new_n432));
  OR3_X1    g0232(.A1(new_n293), .A2(new_n225), .A3(new_n297), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n349), .A3(new_n433), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n434), .A2(G179), .ZN(new_n435));
  INV_X1    g0235(.A(new_n271), .ZN(new_n436));
  OAI21_X1  g0236(.A(G77), .B1(new_n209), .B2(G1), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(G77), .B2(new_n332), .ZN(new_n438));
  INV_X1    g0238(.A(new_n264), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n263), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n438), .B1(new_n443), .B2(new_n267), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n434), .B2(new_n319), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n434), .A2(G200), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n444), .C1(new_n308), .C2(new_n434), .ZN(new_n448));
  AND4_X1   g0248(.A1(new_n422), .A2(new_n427), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n322), .A2(new_n373), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n287), .A2(G244), .A3(new_n383), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT4), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n383), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n453), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n293), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n296), .A2(G1), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n302), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n464), .A2(new_n292), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G257), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n458), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G200), .ZN(new_n468));
  INV_X1    g0268(.A(G33), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n323), .B(new_n332), .C1(G1), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n270), .A2(KEYINPUT82), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT82), .B1(new_n270), .B2(new_n471), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n470), .A2(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g0274(.A1(KEYINPUT81), .A2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT81), .A2(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT6), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n471), .A2(new_n429), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n205), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n483));
  OAI21_X1  g0283(.A(G107), .B1(new_n407), .B2(new_n408), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n474), .B1(new_n485), .B2(new_n267), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n457), .A2(new_n293), .B1(G257), .B2(new_n465), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G190), .A3(new_n461), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n468), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT83), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n468), .A2(new_n486), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  INV_X1    g0292(.A(G179), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n487), .A2(new_n493), .A3(new_n461), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n486), .B1(new_n319), .B2(new_n467), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n490), .A2(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n470), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n441), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n442), .A2(new_n270), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n209), .B(G68), .C1(new_n280), .C2(new_n281), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n263), .B1(new_n475), .B2(new_n476), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(KEYINPUT19), .ZN(new_n502));
  INV_X1    g0302(.A(G87), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n475), .A2(new_n503), .A3(new_n429), .A4(new_n476), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n209), .B1(new_n346), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT84), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(KEYINPUT84), .A3(new_n506), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n267), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n502), .ZN(new_n513));
  INV_X1    g0313(.A(new_n509), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n513), .B(new_n511), .C1(new_n514), .C2(new_n507), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n498), .B(new_n499), .C1(new_n512), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G238), .A2(G1698), .ZN(new_n520));
  INV_X1    g0320(.A(G244), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(new_n522), .B2(new_n287), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n292), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n302), .A2(new_n460), .ZN(new_n525));
  INV_X1    g0325(.A(G250), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n460), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n292), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n493), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n517), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n524), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n302), .A2(new_n460), .B1(new_n527), .B2(new_n292), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(G190), .A4(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(G190), .C1(new_n292), .C2(new_n523), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT86), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n536), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(new_n539), .B1(new_n540), .B2(G200), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n513), .B1(new_n514), .B2(new_n507), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n267), .A3(new_n515), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n497), .A2(G87), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(new_n544), .A3(new_n499), .A4(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT87), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n533), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n533), .B2(new_n546), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n287), .A2(G264), .A3(G1698), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n287), .A2(G257), .A3(new_n383), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n282), .A2(G303), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n293), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n464), .A2(G270), .A3(new_n292), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n461), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G169), .ZN(new_n561));
  INV_X1    g0361(.A(G116), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n270), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n470), .B2(new_n562), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT20), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n455), .A2(new_n209), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n477), .B2(new_n469), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n267), .B1(new_n209), .B2(G116), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n568), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n475), .A2(new_n476), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(G33), .ZN(new_n572));
  OAI211_X1 g0372(.A(KEYINPUT20), .B(new_n570), .C1(new_n572), .C2(new_n566), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n551), .B1(new_n561), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n569), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n497), .A2(G116), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n563), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n578), .A2(KEYINPUT21), .A3(G169), .A4(new_n560), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n558), .B1(new_n293), .B2(new_n555), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n574), .C1(new_n310), .C2(new_n580), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n556), .A2(new_n559), .A3(G179), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  AND4_X1   g0384(.A1(new_n575), .A2(new_n579), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n209), .A2(G107), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n586), .B(KEYINPUT23), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT88), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n518), .B2(G20), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n209), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n287), .A2(new_n209), .A3(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT22), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n287), .A2(new_n594), .A3(new_n209), .A4(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT24), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n591), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n267), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT25), .B1(new_n270), .B2(new_n429), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n429), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n497), .A2(G107), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n464), .A2(G264), .A3(new_n292), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT89), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT89), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n464), .A2(new_n608), .A3(G264), .A4(new_n292), .ZN(new_n609));
  OAI211_X1 g0409(.A(G257), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n610));
  OAI211_X1 g0410(.A(G250), .B(new_n383), .C1(new_n280), .C2(new_n281), .ZN(new_n611));
  INV_X1    g0411(.A(G294), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n611), .C1(new_n469), .C2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n607), .A2(new_n609), .B1(new_n613), .B2(new_n293), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(G179), .A3(new_n461), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(KEYINPUT90), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n293), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n461), .A3(new_n606), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G169), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n615), .B2(KEYINPUT90), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n605), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(G200), .B1(new_n614), .B2(new_n461), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n618), .A2(G190), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n600), .B(new_n604), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n585), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n450), .A2(new_n496), .A3(new_n550), .A4(new_n625), .ZN(G372));
  AND3_X1   g0426(.A1(new_n579), .A2(new_n575), .A3(new_n584), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n538), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(G200), .B2(new_n540), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(new_n544), .A3(new_n499), .A4(new_n545), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n496), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n533), .A2(new_n631), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n495), .A2(new_n494), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT26), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n633), .A2(new_n636), .A3(new_n533), .ZN(new_n637));
  INV_X1    g0437(.A(new_n635), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n550), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n450), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n427), .ZN(new_n643));
  INV_X1    g0443(.A(new_n446), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n372), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n369), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n422), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n315), .B(new_n318), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n321), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n649), .ZN(G369));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n331), .A2(new_n209), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(G213), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n621), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n605), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n621), .A2(new_n624), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n651), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(new_n651), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n627), .A2(new_n657), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n657), .B(KEYINPUT92), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n621), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n665), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n585), .B1(new_n574), .B2(new_n658), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n578), .A2(new_n657), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n627), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n670), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n212), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n504), .A2(G116), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n679), .A2(new_n208), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n221), .B2(new_n679), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n683), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n634), .B2(new_n635), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n633), .A2(new_n688), .A3(new_n533), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT29), .B(new_n658), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n669), .B1(new_n637), .B2(new_n640), .ZN(new_n691));
  XOR2_X1   g0491(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n550), .A2(new_n625), .A3(new_n496), .A4(new_n668), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n580), .A2(new_n614), .A3(new_n530), .A4(G179), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n458), .A2(new_n466), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT30), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n614), .A2(new_n530), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n487), .A4(new_n583), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n580), .A2(new_n530), .A3(G179), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n614), .A2(new_n461), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n467), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n658), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(new_n467), .B1(new_n699), .B2(new_n702), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n668), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n695), .B1(new_n696), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n694), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n686), .B1(new_n717), .B2(G1), .ZN(G364));
  INV_X1    g0518(.A(new_n675), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n269), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n208), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n679), .A2(KEYINPUT95), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT95), .B1(new_n679), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n674), .A2(G330), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n719), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT96), .Z(new_n729));
  NAND2_X1  g0529(.A1(new_n212), .A2(new_n287), .ZN(new_n730));
  INV_X1    g0530(.A(G355), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(G116), .B2(new_n212), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n678), .A2(new_n287), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n296), .B2(new_n221), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n251), .A2(new_n296), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n215), .B1(G20), .B2(new_n319), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n726), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n674), .A2(G20), .A3(new_n739), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n209), .A2(new_n493), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n308), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G326), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(G190), .A3(new_n310), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n287), .B(new_n751), .C1(G322), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(G179), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT99), .Z(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G329), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT97), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n746), .A2(new_n761), .A3(new_n756), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n746), .B2(new_n756), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n754), .B(new_n759), .C1(new_n760), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n747), .A2(G190), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n755), .A2(new_n308), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(G283), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n209), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n770), .B1(new_n612), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n757), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(KEYINPUT32), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n282), .B(new_n778), .C1(G58), .C2(new_n753), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n774), .A2(new_n503), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G50), .B2(new_n748), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n768), .A2(new_n429), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n777), .B2(KEYINPUT32), .ZN(new_n783));
  INV_X1    g0583(.A(new_n764), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G77), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n772), .A2(new_n471), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G68), .B2(new_n766), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT98), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n765), .A2(new_n775), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n744), .B(new_n745), .C1(new_n741), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n729), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  OAI21_X1  g0593(.A(new_n448), .B1(new_n444), .B2(new_n658), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n446), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n644), .A2(new_n658), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n691), .B(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n725), .B1(new_n800), .B2(new_n714), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n714), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n768), .A2(new_n503), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  INV_X1    g0604(.A(new_n766), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(new_n749), .B2(new_n773), .ZN(new_n806));
  INV_X1    g0606(.A(new_n774), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n803), .B(new_n806), .C1(G107), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n758), .A2(G311), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n784), .A2(G116), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n287), .B(new_n787), .C1(G294), .C2(new_n753), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n287), .B1(new_n774), .B2(new_n272), .ZN(new_n813));
  INV_X1    g0613(.A(G58), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n772), .A2(new_n814), .B1(new_n768), .B2(new_n325), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(new_n758), .C2(G132), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G137), .A2(new_n748), .B1(new_n753), .B2(G143), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n260), .B2(new_n805), .C1(new_n391), .C2(new_n764), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n818), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n812), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n824));
  INV_X1    g0624(.A(new_n741), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n823), .B2(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n741), .A2(new_n738), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n725), .B1(new_n226), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n738), .B2(new_n797), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n802), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n720), .A2(new_n208), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  INV_X1    g0635(.A(new_n416), .ZN(new_n836));
  INV_X1    g0636(.A(new_n413), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n406), .A2(new_n267), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n406), .A2(KEYINPUT102), .A3(new_n267), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n387), .A2(new_n388), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n426), .B(KEYINPUT103), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT103), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT16), .B1(new_n409), .B2(new_n412), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n839), .B1(new_n846), .B2(new_n323), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n841), .A3(new_n413), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n843), .B1(new_n848), .B2(new_n416), .ZN(new_n849));
  INV_X1    g0649(.A(new_n426), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n416), .ZN(new_n852));
  INV_X1    g0652(.A(new_n655), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n844), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT105), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n417), .A2(new_n853), .ZN(new_n859));
  AND4_X1   g0659(.A1(new_n418), .A2(new_n426), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n856), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n854), .B1(new_n422), .B2(new_n427), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n860), .B1(new_n855), .B2(KEYINPUT37), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n857), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n835), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n863), .B1(new_n866), .B2(new_n857), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n842), .A2(new_n655), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n426), .B1(new_n842), .B2(new_n843), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n845), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n873), .B2(new_n844), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT105), .B1(new_n874), .B2(new_n860), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT108), .B1(new_n707), .B2(KEYINPUT31), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT108), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n711), .C1(new_n710), .C2(new_n658), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n878), .A2(new_n880), .B1(KEYINPUT31), .B2(new_n707), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n797), .B1(new_n881), .B2(new_n696), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT101), .ZN(new_n883));
  OAI21_X1  g0683(.A(G169), .B1(new_n356), .B2(new_n358), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT14), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n372), .A2(new_n885), .A3(new_n362), .A4(new_n359), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n340), .A2(new_n341), .A3(new_n658), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n369), .A2(new_n889), .A3(new_n372), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n369), .A2(new_n889), .A3(new_n883), .A4(new_n372), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n882), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT40), .B1(new_n877), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AND4_X1   g0695(.A1(KEYINPUT40), .A2(new_n882), .A3(new_n891), .A4(new_n892), .ZN(new_n896));
  INV_X1    g0696(.A(new_n859), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n647), .B2(new_n643), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n418), .A2(new_n426), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n858), .B1(new_n899), .B2(new_n859), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT107), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n860), .A2(KEYINPUT107), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n898), .B(new_n901), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n835), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n876), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n895), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n881), .A2(new_n696), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n450), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n695), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT109), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n907), .C2(new_n909), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n891), .A2(new_n892), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n641), .A2(new_n668), .A3(new_n798), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n796), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n877), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n647), .A2(new_n655), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n869), .B2(new_n875), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT39), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n905), .A2(KEYINPUT39), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT106), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n877), .A2(new_n926), .A3(KEYINPUT39), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n369), .A2(new_n657), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n920), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n450), .B(new_n690), .C1(new_n691), .C2(new_n693), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n649), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n931), .B(new_n933), .Z(new_n934));
  AOI21_X1  g0734(.A(new_n834), .B1(new_n914), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n914), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(G116), .A3(new_n217), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n220), .A2(new_n226), .A3(new_n397), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n325), .A2(G50), .ZN(new_n942));
  OAI211_X1 g0742(.A(G1), .B(new_n269), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n940), .A3(new_n943), .ZN(G367));
  INV_X1    g0744(.A(new_n667), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n496), .B1(new_n486), .B2(new_n668), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n638), .A2(new_n669), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n490), .A2(new_n492), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n951), .B(new_n605), .C1(new_n616), .C2(new_n620), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n669), .B1(new_n952), .B2(new_n635), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n949), .B2(KEYINPUT42), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n544), .A2(new_n499), .A3(new_n545), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n657), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(new_n533), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n533), .A3(new_n631), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n950), .A2(new_n954), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n676), .A2(new_n948), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n965), .B(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n679), .B(KEYINPUT41), .Z(new_n969));
  NOR2_X1   g0769(.A1(new_n665), .A2(new_n666), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n945), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(new_n719), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n716), .ZN(new_n973));
  INV_X1    g0773(.A(new_n948), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n670), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT44), .Z(new_n976));
  INV_X1    g0776(.A(KEYINPUT110), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n676), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n670), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n670), .B2(new_n974), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n981), .A2(new_n983), .B1(new_n977), .B2(new_n676), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n976), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n979), .B1(new_n976), .B2(new_n984), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n969), .B1(new_n988), .B2(new_n717), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n968), .B1(new_n989), .B2(new_n722), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n957), .A2(new_n740), .A3(new_n958), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n805), .A2(new_n391), .B1(new_n768), .B2(new_n226), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n764), .A2(new_n272), .ZN(new_n993));
  INV_X1    g0793(.A(G137), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n287), .B1(new_n757), .B2(new_n994), .C1(new_n752), .C2(new_n260), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n772), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(G68), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n748), .A2(G143), .B1(new_n807), .B2(G58), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n807), .A2(G116), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n282), .B1(new_n752), .B2(new_n773), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G317), .B2(new_n776), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(new_n804), .C2(new_n764), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n766), .A2(G294), .B1(new_n769), .B2(new_n477), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n429), .B2(new_n772), .C1(new_n760), .C2(new_n749), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1000), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n741), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n742), .B1(new_n212), .B2(new_n442), .C1(new_n734), .C2(new_n247), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n991), .A2(new_n726), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n990), .A2(new_n1012), .ZN(G387));
  OAI22_X1  g0813(.A1(new_n730), .A2(new_n680), .B1(G107), .B2(new_n212), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n244), .A2(G45), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT111), .Z(new_n1016));
  AOI211_X1 g0816(.A(G45), .B(new_n681), .C1(G68), .C2(G77), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n264), .A2(G50), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n734), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1014), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n726), .B1(new_n1021), .B2(new_n743), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT112), .Z(new_n1023));
  INV_X1    g0823(.A(G317), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n764), .A2(new_n773), .B1(new_n1024), .B2(new_n752), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT114), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(KEYINPUT114), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n766), .B1(new_n748), .B2(G322), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n997), .A2(G283), .B1(new_n807), .B2(G294), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n282), .B1(new_n757), .B2(new_n750), .C1(new_n562), .C2(new_n768), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n325), .A2(new_n764), .B1(new_n805), .B2(new_n264), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT113), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n287), .B1(new_n757), .B2(new_n260), .C1(new_n752), .C2(new_n272), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n749), .A2(new_n391), .B1(new_n768), .B2(new_n471), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n442), .A2(new_n772), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n774), .A2(new_n226), .ZN(new_n1045));
  OR4_X1    g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1038), .A2(new_n1039), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1023), .B1(new_n741), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT115), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n671), .B2(new_n740), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n972), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n722), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n717), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n973), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n679), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1052), .B1(new_n1053), .B2(new_n1055), .ZN(G393));
  INV_X1    g0856(.A(new_n987), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n721), .B1(new_n1057), .B2(new_n985), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n974), .A2(new_n740), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n742), .B1(new_n212), .B2(new_n571), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n733), .B2(new_n254), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n749), .A2(new_n1024), .B1(new_n760), .B2(new_n752), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT52), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n805), .A2(new_n773), .B1(new_n562), .B2(new_n772), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G283), .B2(new_n807), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n784), .A2(G294), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n287), .B(new_n782), .C1(G322), .C2(new_n776), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n749), .A2(new_n260), .B1(new_n391), .B2(new_n752), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n282), .B(new_n803), .C1(G143), .C2(new_n776), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n997), .A2(G77), .B1(new_n807), .B2(G68), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n784), .A2(new_n439), .B1(G50), .B2(new_n766), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT116), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1068), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n725), .B(new_n1061), .C1(new_n1076), .C2(new_n741), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1058), .B1(new_n1059), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1057), .A2(new_n1054), .A3(new_n985), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n988), .A2(new_n1079), .A3(new_n679), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(G390));
  AOI22_X1  g0881(.A1(new_n691), .A2(new_n795), .B1(new_n644), .B2(new_n658), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n714), .A2(new_n798), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n915), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT117), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n893), .A2(G330), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1085), .A2(KEYINPUT117), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n915), .A2(new_n1084), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n695), .B1(new_n881), .B2(new_n696), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n798), .A2(new_n1092), .B1(new_n891), .B2(new_n892), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n658), .B(new_n795), .C1(new_n687), .C2(new_n689), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n796), .ZN(new_n1095));
  OR3_X1    g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n450), .A2(new_n1092), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n932), .A2(new_n649), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n929), .B1(new_n1082), .B2(new_n915), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n924), .A2(new_n925), .A3(new_n927), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n915), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1095), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n929), .A3(new_n905), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1091), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1087), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1101), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT118), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1101), .B(new_n1112), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1099), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1116), .C1(new_n1117), .C2(new_n1087), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n679), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1117), .B2(new_n1087), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n928), .A2(new_n739), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n287), .B(new_n780), .C1(G116), .C2(new_n753), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n758), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1123), .B1(new_n571), .B2(new_n764), .C1(new_n612), .C2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n997), .A2(G77), .B1(new_n769), .B2(G68), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n429), .B2(new_n805), .C1(new_n804), .C2(new_n749), .ZN(new_n1127));
  INV_X1    g0927(.A(G132), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n287), .B1(new_n752), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G159), .B2(new_n997), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(G125), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1130), .B1(new_n764), .B2(new_n1131), .C1(new_n1124), .C2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n774), .A2(new_n260), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n748), .A2(G128), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n766), .A2(G137), .B1(new_n769), .B2(G50), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1125), .A2(new_n1127), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n741), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n828), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n726), .C1(new_n439), .C2(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1121), .A2(new_n721), .B1(new_n1122), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1120), .A2(new_n1144), .ZN(G378));
  AOI211_X1 g0945(.A(G41), .B(new_n287), .C1(new_n753), .C2(G107), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1146), .A2(new_n998), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n804), .B2(new_n1124), .C1(new_n442), .C2(new_n764), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n805), .A2(new_n471), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n749), .A2(new_n562), .B1(new_n768), .B2(new_n814), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1148), .A2(new_n1045), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(KEYINPUT58), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT58), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n469), .A2(new_n295), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT119), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n272), .C1(G41), .C2(new_n287), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1132), .A2(new_n749), .B1(new_n805), .B2(new_n1128), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G150), .B2(new_n997), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1131), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G128), .A2(new_n753), .B1(new_n807), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1159), .B(new_n1161), .C1(new_n994), .C2(new_n764), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1155), .B1(G124), .B2(new_n776), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n391), .B2(new_n768), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n741), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n726), .C1(G50), .C2(new_n1141), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n313), .A2(new_n655), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n322), .B(new_n1171), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1170), .B1(new_n1174), .B2(new_n738), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n906), .A2(G330), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT121), .B1(new_n1176), .B2(new_n894), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n695), .B1(new_n896), .B2(new_n905), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT121), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n882), .A2(new_n891), .A3(new_n892), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n868), .B2(new_n876), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1178), .B(new_n1179), .C1(KEYINPUT40), .C2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1172), .B(new_n1173), .Z(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1174), .A2(new_n895), .A3(new_n1179), .A4(new_n1178), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1184), .A2(new_n931), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n931), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1175), .B1(new_n1188), .B2(new_n722), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n931), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1184), .A2(new_n931), .A3(new_n1185), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(KEYINPUT57), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1099), .B1(new_n1195), .B2(new_n1116), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n679), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1118), .A2(new_n1100), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1189), .B1(new_n1197), .B2(new_n1199), .ZN(G375));
  NOR2_X1   g1000(.A1(new_n1104), .A2(new_n739), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n562), .A2(new_n805), .B1(new_n749), .B2(new_n612), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1044), .B(new_n1202), .C1(G97), .C2(new_n807), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n282), .B1(new_n768), .B2(new_n226), .C1(new_n804), .C2(new_n752), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G303), .B2(new_n758), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n429), .C2(new_n764), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n749), .A2(new_n1128), .B1(new_n774), .B2(new_n391), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n805), .A2(new_n1131), .B1(new_n272), .B2(new_n772), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n758), .A2(G128), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n784), .A2(G150), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n287), .B1(new_n752), .B2(new_n994), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G58), .B2(new_n769), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1208), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n741), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n726), .C1(G68), .C2(new_n1141), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1201), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1097), .B2(new_n722), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1116), .A2(new_n969), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1090), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G387), .A2(new_n1230), .A3(G378), .A4(G375), .ZN(G407));
  AOI21_X1  g1031(.A(new_n1143), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n656), .A2(G213), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G407), .B(G213), .C1(G375), .C2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n1099), .A4(new_n1096), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1239), .A2(new_n679), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1225), .B1(new_n1116), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1243), .A2(G384), .A3(new_n1222), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G384), .B1(new_n1243), .B2(new_n1222), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(G2897), .A3(new_n1234), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1234), .A2(G2897), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1251), .B2(new_n1248), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT57), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1196), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1188), .A2(new_n1198), .A3(KEYINPUT57), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n679), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(G378), .A3(new_n1189), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n969), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1188), .A2(new_n1198), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1189), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1232), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1234), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1238), .B1(new_n1252), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n990), .B2(new_n1012), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n990), .A2(G390), .A3(new_n1012), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n792), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1266), .A2(new_n1270), .A3(new_n1269), .A4(new_n1267), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1264), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1262), .B1(G375), .B2(new_n1232), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1233), .A3(new_n1246), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT124), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1263), .A2(new_n1279), .A3(new_n1246), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1246), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1275), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1276), .A2(KEYINPUT62), .A3(new_n1233), .A4(new_n1246), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT127), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1263), .A2(new_n1287), .A3(KEYINPUT62), .A4(new_n1246), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1278), .A2(new_n1280), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1264), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1274), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1284), .B1(new_n1292), .B2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1232), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1258), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1246), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1296), .B(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1293), .B(new_n1298), .ZN(G402));
endmodule


