//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n224), .A2(G50), .A3(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n207), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n212), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT80), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n253), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G116), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n257), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n228), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n206), .B2(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G283), .ZN(new_n265));
  INV_X1    g0065(.A(G97), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n265), .B(new_n207), .C1(G33), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT79), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(G20), .B1(new_n269), .B2(G97), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT79), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(new_n265), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n260), .A2(new_n228), .B1(G20), .B2(new_n255), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n273), .A2(KEYINPUT20), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT20), .B1(new_n273), .B2(new_n274), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n258), .B(new_n264), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n269), .ZN(new_n282));
  INV_X1    g0082(.A(G303), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G257), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G264), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G1698), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n280), .B(new_n285), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT5), .B(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n293), .A2(G274), .A3(new_n279), .A4(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT5), .A2(G41), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT5), .A2(G41), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G270), .A3(new_n279), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n292), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n250), .B1(new_n277), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT21), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n264), .A2(new_n258), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n273), .A2(new_n274), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n273), .A2(KEYINPUT20), .A3(new_n274), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND4_X1   g0111(.A1(G179), .A2(new_n292), .A3(new_n296), .A4(new_n300), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n304), .A2(new_n305), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT80), .B1(new_n311), .B2(new_n302), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(KEYINPUT21), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n301), .A2(G200), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n301), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n277), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n314), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n207), .A2(G33), .ZN(new_n323));
  INV_X1    g0123(.A(G150), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G20), .A2(G33), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n322), .A2(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G50), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n207), .B1(new_n223), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n261), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n256), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n261), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n206), .A2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(G50), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n330), .B(new_n334), .C1(G50), .C2(new_n256), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT70), .ZN(new_n338));
  INV_X1    g0138(.A(G41), .ZN(new_n339));
  AOI21_X1  g0139(.A(G1), .B1(new_n339), .B2(new_n294), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(new_n279), .A3(G274), .ZN(new_n341));
  INV_X1    g0141(.A(G226), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n279), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(KEYINPUT67), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n282), .A2(new_n284), .ZN(new_n347));
  INV_X1    g0147(.A(G1698), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(G222), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(G223), .A3(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G77), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(new_n347), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n280), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n345), .A2(KEYINPUT67), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n346), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(new_n318), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n335), .A2(new_n336), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G200), .B2(new_n355), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n338), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT10), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n335), .C1(G179), .C2(new_n355), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n347), .A2(G232), .A3(new_n348), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n347), .A2(G238), .A3(G1698), .ZN(new_n365));
  INV_X1    g0165(.A(G107), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n347), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n280), .ZN(new_n368));
  INV_X1    g0168(.A(new_n341), .ZN(new_n369));
  INV_X1    g0169(.A(new_n344), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(G244), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n318), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n261), .B1(new_n254), .B2(new_n257), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(G77), .A3(new_n333), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G20), .A2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n376), .B1(new_n377), .B2(new_n323), .C1(new_n326), .C2(new_n322), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n261), .ZN(new_n379));
  INV_X1    g0179(.A(new_n259), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n380), .A2(KEYINPUT69), .A3(new_n351), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT69), .B1(new_n380), .B2(new_n351), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n375), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n372), .A2(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n372), .A2(new_n361), .ZN(new_n387));
  INV_X1    g0187(.A(G179), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n368), .A2(new_n388), .A3(new_n371), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n360), .A2(new_n363), .A3(new_n386), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n202), .A2(G20), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n392), .B1(new_n323), .B2(new_n351), .C1(new_n326), .C2(new_n328), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n261), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT11), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n374), .A2(G68), .A3(new_n333), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n392), .A2(KEYINPUT12), .A3(G1), .A4(new_n251), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n380), .A2(new_n202), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(KEYINPUT12), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT13), .ZN(new_n404));
  OAI211_X1 g0204(.A(G226), .B(new_n348), .C1(new_n289), .C2(new_n290), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n347), .A2(KEYINPUT71), .A3(G226), .A4(new_n348), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n347), .A2(G232), .A3(G1698), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n280), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n341), .B1(new_n214), .B2(new_n344), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n404), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI211_X1 g0215(.A(KEYINPUT13), .B(new_n413), .C1(new_n411), .C2(new_n280), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n403), .B(G169), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n414), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n388), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n403), .B1(new_n421), .B2(G169), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n402), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n415), .A2(new_n416), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G190), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n415), .B2(new_n416), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n401), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G58), .A2(G68), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n207), .B1(new_n203), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n325), .A2(G159), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n431), .ZN(new_n436));
  OAI21_X1  g0236(.A(G20), .B1(new_n436), .B2(new_n223), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT73), .A3(new_n433), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT72), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n282), .A2(new_n207), .A3(new_n284), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT7), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n284), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(new_n446), .B2(G68), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT72), .B(new_n202), .C1(new_n444), .C2(new_n445), .ZN(new_n448));
  OAI211_X1 g0248(.A(KEYINPUT16), .B(new_n440), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT16), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n202), .B1(new_n444), .B2(new_n445), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n439), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n261), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n332), .ZN(new_n454));
  INV_X1    g0254(.A(new_n322), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n333), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n454), .A2(new_n456), .B1(new_n256), .B2(new_n455), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n279), .A2(G232), .A3(new_n343), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n341), .A2(new_n460), .A3(KEYINPUT74), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT74), .B1(new_n341), .B2(new_n460), .ZN(new_n462));
  OR2_X1    g0262(.A1(G223), .A2(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n342), .A2(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n464), .C1(new_n289), .C2(new_n290), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G87), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n279), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n461), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G179), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n341), .A2(new_n460), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT74), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n280), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n341), .A2(new_n460), .A3(KEYINPUT74), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G169), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n459), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT18), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n318), .ZN(new_n481));
  OAI211_X1 g0281(.A(KEYINPUT75), .B(new_n481), .C1(new_n468), .C2(G200), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G200), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT75), .B1(new_n485), .B2(new_n481), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n453), .B(new_n458), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT17), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT18), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n459), .A2(new_n478), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT75), .ZN(new_n492));
  INV_X1    g0292(.A(new_n481), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n462), .A2(new_n467), .ZN(new_n494));
  AOI21_X1  g0294(.A(G200), .B1(new_n494), .B2(new_n475), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n482), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT17), .A3(new_n453), .A4(new_n458), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n480), .A2(new_n489), .A3(new_n491), .A4(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n391), .A2(new_n429), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n332), .B1(G1), .B2(new_n269), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n366), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n331), .A2(new_n366), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT25), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n207), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT22), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT22), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n347), .A2(new_n509), .A3(new_n207), .A4(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G20), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT23), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n207), .B2(G107), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n366), .A2(KEYINPUT23), .A3(G20), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n511), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n506), .B1(new_n522), .B2(new_n261), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n279), .A2(G274), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(new_n299), .ZN(new_n525));
  INV_X1    g0325(.A(G257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G1698), .ZN(new_n527));
  OAI221_X1 g0327(.A(new_n527), .B1(G250), .B2(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G294), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n525), .B1(new_n530), .B2(new_n280), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n299), .A2(G264), .A3(new_n279), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n361), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n299), .A2(new_n535), .A3(G264), .A4(new_n279), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n279), .B1(new_n528), .B2(new_n529), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n537), .A2(new_n296), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n533), .B1(new_n540), .B2(G179), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n501), .B1(new_n523), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n521), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n520), .B1(new_n511), .B2(new_n517), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n261), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n503), .A2(new_n505), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n537), .A2(new_n296), .A3(new_n539), .ZN(new_n548));
  INV_X1    g0348(.A(new_n532), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n538), .A2(new_n549), .A3(new_n525), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n548), .A2(new_n388), .B1(new_n550), .B2(new_n361), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n551), .A3(KEYINPUT82), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G250), .A2(G1698), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT4), .A2(G244), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(G1698), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n347), .A2(new_n556), .B1(G33), .B2(G283), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(new_n348), .C1(new_n289), .C2(new_n290), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n279), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n299), .A2(new_n279), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n296), .B1(new_n562), .B2(new_n526), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n388), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n361), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n446), .A2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n366), .A2(KEYINPUT6), .A3(G97), .ZN(new_n568));
  AND2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n571), .B2(KEYINPUT6), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G20), .B1(G77), .B2(new_n325), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n262), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n331), .A2(new_n266), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n502), .B2(new_n266), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n565), .B(new_n566), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n567), .A2(new_n573), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n576), .B1(new_n578), .B2(new_n261), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n564), .A2(G190), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n561), .B2(new_n563), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n548), .A2(new_n484), .B1(new_n550), .B2(new_n318), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n577), .B(new_n582), .C1(new_n547), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n215), .A2(new_n266), .A3(new_n366), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT77), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(new_n215), .A3(new_n266), .A4(new_n366), .ZN(new_n588));
  NAND3_X1  g0388(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n586), .A2(new_n588), .B1(new_n207), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n207), .B(G68), .C1(new_n289), .C2(new_n290), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n323), .B2(new_n266), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n261), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n380), .A2(new_n377), .ZN(new_n596));
  INV_X1    g0396(.A(new_n377), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n332), .B(new_n597), .C1(G1), .C2(new_n269), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT78), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n595), .A2(new_n601), .A3(new_n596), .A4(new_n598), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n295), .A2(new_n216), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n279), .ZN(new_n604));
  INV_X1    g0404(.A(new_n295), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n524), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT76), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n347), .A2(KEYINPUT76), .A3(G244), .A4(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n347), .A2(G238), .A3(new_n348), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n512), .A4(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n606), .B1(new_n612), .B2(new_n280), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(new_n361), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n388), .B(new_n606), .C1(new_n612), .C2(new_n280), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n600), .B(new_n602), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n595), .A2(new_n596), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n502), .A2(new_n215), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(G190), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n484), .C2(new_n613), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n584), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n321), .A2(new_n500), .A3(new_n553), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g0424(.A(new_n624), .B(KEYINPUT83), .Z(G372));
  AND2_X1   g0425(.A1(new_n480), .A2(new_n491), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT14), .B1(new_n425), .B2(new_n361), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n417), .C1(new_n388), .C2(new_n421), .ZN(new_n628));
  INV_X1    g0428(.A(new_n390), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n628), .A2(new_n402), .B1(new_n428), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n489), .A2(new_n498), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n360), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n363), .ZN(new_n634));
  INV_X1    g0434(.A(new_n500), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n599), .B1(new_n614), .B2(new_n615), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n621), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(new_n566), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n561), .A2(new_n563), .A3(G179), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n579), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n616), .A2(new_n642), .A3(new_n621), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n636), .B(KEYINPUT84), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n584), .A2(new_n637), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n311), .A2(new_n313), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n315), .B2(KEYINPUT21), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n304), .A2(new_n305), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n547), .A2(new_n551), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n634), .B1(new_n635), .B2(new_n657), .ZN(G369));
  XNOR2_X1  g0458(.A(KEYINPUT86), .B(G330), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n252), .A2(new_n207), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT85), .Z(new_n661));
  INV_X1    g0461(.A(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G213), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n321), .B1(new_n311), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n277), .B(new_n667), .C1(new_n314), .C2(new_n316), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n659), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n547), .A2(new_n583), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n547), .B2(new_n667), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n553), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n547), .A2(new_n667), .A3(new_n551), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n668), .A2(new_n547), .A3(new_n551), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n667), .B1(new_n651), .B2(new_n652), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n553), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n210), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT87), .B1(new_n682), .B2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n682), .A2(KEYINPUT87), .A3(G41), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n586), .A2(new_n255), .A3(new_n588), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n226), .B2(new_n687), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n649), .A2(new_n654), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n693), .B(new_n668), .C1(new_n694), .C2(new_n647), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n644), .A2(new_n639), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n638), .A2(KEYINPUT26), .A3(new_n642), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n644), .A2(KEYINPUT90), .A3(new_n639), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n542), .A2(new_n652), .A3(new_n651), .A4(new_n552), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n584), .A2(new_n637), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT91), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n703), .B2(new_n704), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n702), .B(new_n646), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n668), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n696), .B1(new_n709), .B2(KEYINPUT29), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n538), .B1(new_n534), .B2(new_n536), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n564), .A2(new_n711), .A3(new_n312), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT88), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT30), .A4(new_n613), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n613), .A2(new_n564), .A3(new_n711), .A4(new_n312), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT88), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n613), .ZN(new_n719));
  INV_X1    g0519(.A(new_n564), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n301), .A2(new_n388), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n548), .A4(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT89), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n715), .B2(new_n716), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n715), .A2(new_n723), .A3(new_n716), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n718), .A2(new_n722), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n667), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n553), .A2(new_n321), .A3(new_n623), .A4(new_n668), .ZN(new_n731));
  INV_X1    g0531(.A(new_n722), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n714), .B2(new_n717), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n715), .A2(new_n716), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n659), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n710), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n692), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n251), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n206), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n686), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n671), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n669), .A2(new_n659), .A3(new_n670), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n669), .A2(new_n670), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n745), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n682), .A2(new_n291), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G355), .B1(new_n255), .B2(new_n682), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n682), .A2(new_n347), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G45), .B2(new_n226), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n248), .A2(new_n294), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n228), .B1(G20), .B2(new_n361), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n751), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n753), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT92), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(KEYINPUT92), .ZN(new_n764));
  INV_X1    g0564(.A(new_n760), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n318), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n207), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n207), .A2(new_n388), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n767), .A2(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n318), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(G326), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(G190), .A3(new_n484), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n291), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n770), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(G329), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n774), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n781), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n781), .A2(new_n318), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(G303), .B1(new_n793), .B2(G283), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n777), .A2(new_n784), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n775), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT32), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n782), .A2(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n796), .A2(new_n328), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G68), .B2(new_n785), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n347), .B1(new_n771), .B2(new_n351), .ZN(new_n802));
  INV_X1    g0602(.A(new_n778), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G58), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n767), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G97), .B1(new_n791), .B2(G87), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n797), .A2(new_n799), .B1(new_n793), .B2(G107), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n801), .A2(new_n804), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n765), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n764), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n752), .A2(new_n763), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n748), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  AOI21_X1  g0613(.A(new_n667), .B1(new_n648), .B2(new_n655), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n390), .A2(KEYINPUT94), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT94), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n387), .A2(new_n383), .A3(new_n816), .A4(new_n389), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n818), .A2(new_n386), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n667), .A2(new_n383), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n386), .A2(new_n815), .A3(new_n821), .A4(new_n817), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n629), .A2(new_n667), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n820), .B1(new_n814), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n745), .B1(new_n825), .B2(new_n739), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n739), .B2(new_n825), .ZN(new_n827));
  INV_X1    g0627(.A(new_n771), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n803), .A2(G143), .B1(new_n828), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(new_n785), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n796), .B2(new_n830), .C1(new_n324), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n792), .A2(new_n202), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n291), .B(new_n836), .C1(G132), .C2(new_n783), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n805), .A2(G58), .B1(new_n791), .B2(G50), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n796), .A2(new_n283), .B1(new_n790), .B2(new_n366), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G87), .B2(new_n793), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n347), .B1(new_n803), .B2(G294), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G116), .A2(new_n828), .B1(new_n783), .B2(G311), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G97), .A2(new_n805), .B1(new_n785), .B2(G283), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n765), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n760), .A2(new_n749), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n753), .B(new_n846), .C1(new_n351), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n824), .B2(new_n750), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n827), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  OR2_X1    g0651(.A1(new_n572), .A2(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n572), .A2(KEYINPUT35), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(G116), .A3(new_n229), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n855));
  XNOR2_X1  g0655(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n227), .A2(G77), .A3(new_n431), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n328), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n206), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT7), .B1(new_n291), .B2(new_n207), .ZN(new_n861));
  INV_X1    g0661(.A(new_n445), .ZN(new_n862));
  OAI21_X1  g0662(.A(G68), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT72), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n451), .A2(new_n441), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n439), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n262), .B1(new_n866), .B2(KEYINPUT16), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n440), .B1(new_n447), .B2(new_n448), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n450), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n457), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n664), .A2(new_n666), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n487), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n469), .A2(new_n477), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n459), .A2(new_n871), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n479), .A2(new_n877), .A3(new_n487), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n870), .A2(new_n872), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n499), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n880), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n428), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n402), .B(new_n667), .C1(new_n628), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n402), .A2(new_n667), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n424), .A2(new_n428), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n820), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n818), .A2(new_n667), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n887), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n877), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n499), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n479), .A2(new_n877), .A3(new_n487), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n879), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n885), .B(new_n886), .C1(KEYINPUT96), .C2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n901), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT96), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(KEYINPUT39), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n902), .A2(KEYINPUT39), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n628), .A2(new_n402), .A3(new_n668), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n895), .B1(new_n626), .B2(new_n871), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n634), .B1(new_n710), .B2(new_n635), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n909), .B(new_n910), .Z(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n880), .B2(new_n882), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n903), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n730), .A2(new_n915), .A3(new_n731), .ZN(new_n916));
  INV_X1    g0716(.A(new_n824), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n889), .B2(new_n891), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n499), .A2(new_n896), .B1(new_n899), .B2(new_n879), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n886), .B1(KEYINPUT38), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n916), .A2(new_n918), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n912), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n500), .A2(new_n916), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n659), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n911), .A2(new_n928), .B1(new_n206), .B2(new_n742), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n911), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n860), .B1(new_n929), .B2(new_n930), .ZN(G367));
  INV_X1    g0731(.A(new_n619), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n667), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n646), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n638), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n936), .A2(G20), .A3(new_n750), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n756), .A2(new_n235), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(new_n761), .C1(new_n210), .C2(new_n377), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n831), .A2(new_n768), .B1(new_n792), .B2(new_n266), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n796), .A2(new_n772), .B1(new_n366), .B2(new_n767), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(G283), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n291), .B1(new_n771), .B2(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n778), .A2(new_n283), .B1(new_n782), .B2(new_n786), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n790), .A2(new_n255), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n944), .B(new_n945), .C1(KEYINPUT46), .C2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n942), .B(new_n947), .C1(KEYINPUT46), .C2(new_n946), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n831), .A2(new_n798), .B1(new_n202), .B2(new_n767), .ZN(new_n949));
  INV_X1    g0749(.A(G143), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n796), .A2(new_n950), .B1(new_n790), .B2(new_n201), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n778), .A2(new_n324), .B1(new_n771), .B2(new_n328), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G137), .B2(new_n783), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n291), .B1(new_n793), .B2(G77), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT105), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n952), .A2(new_n954), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n948), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  OAI211_X1 g0760(.A(new_n745), .B(new_n939), .C1(new_n960), .C2(new_n765), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n937), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT100), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n577), .B(new_n582), .C1(new_n668), .C2(new_n579), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n642), .A2(new_n667), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n967), .A2(new_n553), .A3(new_n673), .A4(new_n679), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n577), .B1(new_n553), .B2(new_n965), .ZN(new_n969));
  AOI22_X1  g0769(.A1(KEYINPUT42), .A2(new_n968), .B1(new_n969), .B2(new_n668), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n934), .A2(new_n975), .A3(new_n935), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT97), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n964), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n972), .A2(new_n973), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(KEYINPUT100), .A3(new_n978), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT99), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT98), .B1(new_n981), .B2(new_n978), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT98), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n986), .A3(new_n974), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n983), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n985), .A2(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n980), .A2(new_n982), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT99), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n967), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n989), .A2(new_n992), .B1(new_n677), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n984), .B1(new_n983), .B2(new_n988), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n677), .A2(new_n993), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n990), .A2(KEYINPUT99), .A3(new_n991), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n680), .A2(new_n678), .A3(new_n967), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT101), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT101), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n680), .A2(new_n678), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n993), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT103), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(KEYINPUT44), .A3(new_n993), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(KEYINPUT103), .A3(new_n1013), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1005), .A2(new_n1006), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n677), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1014), .A2(new_n1011), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1018), .A2(new_n677), .A3(new_n1006), .A4(new_n1005), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT104), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n680), .B1(new_n676), .B2(new_n679), .C1(new_n671), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n671), .A2(new_n1021), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n740), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n740), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n686), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n744), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n963), .B1(new_n999), .B2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n1025), .A2(new_n686), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1024), .A2(new_n740), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n674), .A2(new_n675), .A3(new_n751), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G311), .A2(new_n785), .B1(new_n775), .B2(G322), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT108), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(KEYINPUT108), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n803), .A2(G317), .B1(new_n828), .B2(G303), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n805), .A2(G283), .B1(new_n791), .B2(G294), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n792), .A2(new_n255), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n347), .B(new_n1048), .C1(G326), .C2(new_n783), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n771), .A2(new_n202), .B1(new_n782), .B2(new_n324), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n291), .B(new_n1051), .C1(G50), .C2(new_n803), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n791), .A2(G77), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n597), .A2(new_n805), .B1(new_n785), .B2(new_n455), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n775), .A2(G159), .B1(new_n793), .B2(G97), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n765), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n689), .B(new_n294), .C1(new_n202), .C2(new_n351), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT106), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n322), .A2(G50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT50), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1058), .B2(KEYINPUT106), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n756), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT107), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n294), .C2(new_n240), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n754), .A2(new_n688), .B1(new_n366), .B2(new_n682), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n753), .B(new_n1057), .C1(new_n761), .C2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1024), .A2(new_n744), .B1(new_n1034), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1033), .A2(new_n1071), .ZN(G393));
  NOR2_X1   g0872(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1073), .A2(new_n687), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT109), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT109), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1025), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n993), .A2(new_n751), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n245), .A2(new_n682), .A3(new_n347), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n761), .B1(new_n266), .B2(new_n210), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n796), .A2(new_n324), .B1(new_n798), .B2(new_n778), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n831), .A2(new_n328), .B1(new_n792), .B2(new_n215), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n347), .B1(new_n782), .B2(new_n950), .C1(new_n322), .C2(new_n771), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n767), .A2(new_n351), .B1(new_n790), .B2(new_n202), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n796), .A2(new_n786), .B1(new_n772), .B2(new_n778), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n831), .A2(new_n283), .B1(new_n255), .B2(new_n767), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n291), .B1(new_n782), .B2(new_n779), .C1(new_n768), .C2(new_n771), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n366), .A2(new_n792), .B1(new_n790), .B2(new_n943), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1083), .A2(new_n1087), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n745), .B1(new_n1080), .B2(new_n1081), .C1(new_n1094), .C2(new_n765), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT111), .Z(new_n1096));
  AOI22_X1  g0896(.A1(new_n1074), .A2(new_n1078), .B1(new_n1079), .B2(new_n1096), .ZN(new_n1097));
  OR3_X1    g0897(.A1(new_n1076), .A2(KEYINPUT110), .A3(new_n1077), .ZN(new_n1098));
  OAI21_X1  g0898(.A(KEYINPUT110), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n744), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(G390));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n778), .A2(new_n1102), .B1(new_n782), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n291), .B(new_n1104), .C1(new_n828), .C2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n790), .A2(new_n324), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G159), .A2(new_n805), .B1(new_n785), .B2(G137), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n775), .A2(G128), .B1(new_n793), .B2(G50), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n291), .B1(new_n790), .B2(new_n215), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT113), .Z(new_n1114));
  OAI22_X1  g0914(.A1(new_n771), .A2(new_n266), .B1(new_n782), .B2(new_n768), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G116), .B2(new_n803), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n836), .B1(G77), .B2(new_n805), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G107), .A2(new_n785), .B1(new_n775), .B2(G283), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n765), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n753), .B(new_n1120), .C1(new_n322), .C2(new_n847), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n907), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n750), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n894), .B1(new_n814), .B2(new_n819), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n892), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n908), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n904), .A2(new_n906), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1124), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n708), .A2(new_n668), .A3(new_n819), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n894), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n892), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n922), .A2(new_n908), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n737), .A2(new_n738), .A3(new_n824), .A4(new_n892), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n916), .A2(new_n918), .A3(G330), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(KEYINPUT112), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1129), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n907), .A2(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n916), .A2(G330), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(KEYINPUT112), .A3(new_n918), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1140), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1123), .B1(new_n1145), .B2(new_n743), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n500), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(new_n634), .C1(new_n710), .C2(new_n635), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n737), .A2(new_n738), .A3(new_n824), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1126), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1138), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n893), .B2(new_n894), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1126), .B1(new_n1142), .B2(new_n917), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(new_n1131), .A3(new_n1130), .A4(new_n1136), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n1140), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n687), .B1(new_n1145), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1146), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(G378));
  OAI211_X1 g0960(.A(KEYINPUT117), .B(G330), .C1(new_n920), .C2(new_n924), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n360), .A2(new_n363), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n360), .A2(new_n363), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n871), .A2(new_n335), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT115), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1167), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1161), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT40), .B1(new_n904), .B2(new_n919), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n887), .A2(new_n912), .A3(new_n923), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT117), .B1(new_n1175), .B2(G330), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g0977(.A(KEYINPUT117), .B(new_n1171), .C1(new_n1175), .C2(G330), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n909), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1148), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1156), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT117), .ZN(new_n1182));
  INV_X1    g0982(.A(G330), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n925), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n1161), .A3(new_n1171), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n909), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1179), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1179), .A2(new_n1181), .A3(new_n1188), .A4(KEYINPUT57), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n686), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1179), .A2(new_n744), .A3(new_n1188), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1171), .A2(new_n749), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n796), .A2(new_n255), .B1(new_n792), .B2(new_n201), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G97), .B2(new_n785), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n291), .A2(new_n339), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G283), .B2(new_n783), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n803), .A2(G107), .B1(new_n828), .B2(new_n597), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n805), .A2(G68), .B1(new_n791), .B2(G77), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G50), .B1(new_n269), .B2(new_n339), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1202), .A2(new_n1203), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n785), .A2(G132), .B1(new_n828), .B2(G137), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT114), .ZN(new_n1207));
  INV_X1    g1007(.A(G128), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n767), .A2(new_n324), .B1(new_n778), .B2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n796), .A2(new_n1103), .B1(new_n790), .B2(new_n1105), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n793), .A2(G159), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1205), .B1(new_n1203), .B2(new_n1202), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n760), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n753), .B1(new_n328), .B2(new_n847), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1195), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT116), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1194), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1193), .A2(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n744), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1126), .A2(new_n749), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT118), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n255), .A2(new_n831), .B1(new_n796), .B2(new_n768), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G97), .B2(new_n791), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n793), .A2(G77), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n805), .A2(new_n597), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n778), .A2(new_n943), .B1(new_n771), .B2(new_n366), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n347), .B(new_n1234), .C1(G303), .C2(new_n783), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n347), .B1(new_n792), .B2(new_n201), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT119), .Z(new_n1238));
  OAI22_X1  g1038(.A1(new_n790), .A2(new_n798), .B1(new_n782), .B2(new_n1208), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT120), .Z(new_n1240));
  OAI22_X1  g1040(.A1(new_n778), .A2(new_n830), .B1(new_n771), .B2(new_n324), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G132), .B2(new_n775), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G50), .A2(new_n805), .B1(new_n785), .B2(new_n1106), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1236), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n760), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n847), .A2(new_n202), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1229), .A2(new_n745), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1227), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1155), .A2(new_n1027), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1226), .A2(new_n1180), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1252), .B2(new_n1253), .ZN(G381));
  NOR3_X1   g1054(.A1(G390), .A2(G387), .A3(G381), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1033), .A2(new_n1071), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n812), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT121), .B1(new_n1258), .B2(new_n850), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT121), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1257), .A2(new_n1260), .A3(G384), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1255), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT122), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G378), .B1(G375), .B2(KEYINPUT123), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(KEYINPUT123), .B2(G375), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1263), .A2(new_n1265), .ZN(G407));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G343), .C2(new_n1265), .ZN(G409));
  INV_X1    g1067(.A(new_n998), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1029), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G390), .A2(new_n1272), .A3(new_n963), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G387), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1257), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n962), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT126), .B1(new_n1279), .B2(G390), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1275), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1273), .A2(new_n1274), .A3(KEYINPUT126), .A4(new_n1277), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1281), .A2(KEYINPUT127), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT127), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n665), .A2(G213), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n687), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1159), .B(new_n1223), .C1(new_n1288), .C2(new_n1192), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1194), .B(new_n1221), .C1(new_n1189), .C2(new_n1027), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1159), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1287), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1152), .A2(new_n1148), .A3(KEYINPUT60), .A4(new_n1154), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n686), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1157), .A2(KEYINPUT60), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1253), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1298), .A2(new_n850), .A3(new_n1249), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n850), .B1(new_n1298), .B2(new_n1249), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(G2897), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1287), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1287), .A2(new_n1303), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1300), .A2(new_n1301), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT62), .B1(new_n1293), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1302), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1287), .B(new_n1309), .C1(new_n1289), .C2(new_n1292), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1286), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(KEYINPUT124), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1193), .A2(G378), .A3(new_n1224), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1291), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT124), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n1287), .A4(new_n1309), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT62), .B1(new_n1313), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1285), .B1(new_n1312), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1313), .A2(new_n1320), .A3(new_n1317), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT125), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1304), .A2(new_n1324), .A3(new_n1306), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1293), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1321), .A2(new_n1322), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1159), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1314), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1309), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1285), .B(new_n1332), .ZN(G402));
endmodule


