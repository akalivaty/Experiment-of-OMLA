//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G146), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n194), .B1(new_n193), .B2(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G237), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G953), .ZN(new_n201));
  INV_X1    g015(.A(G953), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT71), .ZN(new_n203));
  OAI211_X1 g017(.A(G214), .B(new_n199), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(KEYINPUT71), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(G953), .ZN(new_n209));
  AOI21_X1  g023(.A(G237), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(G143), .A3(G214), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT18), .A2(G131), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n206), .B(new_n211), .C1(KEYINPUT87), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n215), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n198), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  INV_X1    g034(.A(new_n191), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT19), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT19), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n191), .A2(KEYINPUT90), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n227));
  OR3_X1    g041(.A1(new_n191), .A2(KEYINPUT79), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT79), .B1(new_n191), .B2(new_n227), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n187), .A3(G125), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n229), .A3(G146), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n206), .B2(new_n211), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n206), .A2(new_n233), .A3(new_n211), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT91), .B1(new_n219), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G113), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n236), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n231), .B(new_n226), .C1(new_n243), .C2(new_n234), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n214), .A2(new_n216), .B1(new_n215), .B2(new_n212), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n244), .B(new_n245), .C1(new_n246), .C2(new_n198), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n238), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n235), .A2(new_n249), .A3(new_n236), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT92), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n228), .A2(new_n230), .A3(new_n229), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n220), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n231), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT92), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n235), .A2(new_n257), .A3(new_n249), .A4(new_n236), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n255), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n219), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n241), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G475), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT20), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT93), .ZN(new_n267));
  AOI21_X1  g081(.A(G475), .B1(new_n248), .B2(new_n261), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  AND4_X1   g085(.A1(new_n269), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT93), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n259), .A2(new_n260), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n242), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n261), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n263), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n271), .A2(new_n273), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT99), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT69), .B(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G143), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT95), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G134), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n205), .A2(G128), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n283), .B(KEYINPUT95), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n287), .B(KEYINPUT13), .Z(new_n291));
  OAI21_X1  g105(.A(G134), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT96), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT96), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(G134), .C1(new_n290), .C2(new_n291), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n296));
  INV_X1    g110(.A(G122), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(G116), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT94), .A3(G122), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n298), .A2(new_n300), .B1(G116), .B2(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(G107), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n289), .A2(new_n293), .A3(new_n295), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(G116), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n305), .B2(KEYINPUT14), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n301), .B(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n288), .B2(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT9), .B(G234), .Z(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n304), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n304), .B2(new_n309), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n264), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G478), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI221_X1 g134(.A(new_n264), .B1(KEYINPUT15), .B2(new_n318), .C1(new_n315), .C2(new_n316), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n202), .A2(G952), .ZN(new_n323));
  NAND2_X1  g137(.A1(G234), .A2(G237), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n325), .B(KEYINPUT97), .Z(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n208), .A2(new_n209), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(G902), .A3(new_n324), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT21), .B(G898), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT98), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n322), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n280), .A2(new_n281), .A3(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n322), .A2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT99), .B1(new_n279), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n282), .A2(G119), .ZN(new_n341));
  INV_X1    g155(.A(G128), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(G119), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT77), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT24), .B(G110), .Z(new_n345));
  OR2_X1    g159(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n347));
  INV_X1    g161(.A(G119), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(G128), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n350));
  OAI221_X1 g164(.A(new_n349), .B1(G119), .B2(new_n342), .C1(new_n341), .C2(new_n350), .ZN(new_n351));
  OAI22_X1  g165(.A1(new_n344), .A2(new_n345), .B1(G110), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n231), .A3(new_n193), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n344), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(G110), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n254), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n328), .A2(G221), .A3(G234), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n358), .B(KEYINPUT22), .Z(new_n359));
  INV_X1    g173(.A(G137), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n356), .A3(new_n361), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n264), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n365), .B2(G902), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(G217), .A2(G902), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n312), .B2(G234), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT76), .Z(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G902), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n370), .A2(new_n373), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G472), .A2(G902), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n205), .A2(G146), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n220), .A2(G143), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G128), .ZN(new_n382));
  AND2_X1   g196(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n383));
  NOR2_X1   g197(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G143), .B(G146), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT68), .A4(G128), .ZN(new_n389));
  OR2_X1    g203(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n381), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(KEYINPUT69), .A2(G128), .ZN(new_n393));
  NOR2_X1   g207(.A1(KEYINPUT69), .A2(G128), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n220), .A2(KEYINPUT64), .A3(G143), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT64), .B1(new_n220), .B2(G143), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n380), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n386), .A2(new_n389), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n286), .A2(G137), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n360), .A2(G134), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G131), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT66), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT11), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n286), .B2(G137), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n360), .A2(KEYINPUT11), .A3(G134), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n233), .A4(new_n401), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n404), .A2(KEYINPUT66), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n400), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n401), .A3(new_n408), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G131), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n409), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT0), .B(G128), .Z(new_n417));
  AND3_X1   g231(.A1(new_n380), .A2(new_n381), .A3(G128), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n399), .A2(new_n417), .B1(new_n418), .B2(KEYINPUT0), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(KEYINPUT65), .A3(G131), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n378), .B1(new_n412), .B2(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT2), .B(G113), .Z(new_n423));
  NAND2_X1  g237(.A1(new_n348), .A2(G116), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n299), .A2(G119), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT2), .B(G113), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n386), .A2(new_n389), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n396), .A2(new_n399), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n405), .A2(new_n409), .ZN(new_n434));
  INV_X1    g248(.A(new_n411), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n422), .A2(new_n430), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n430), .B(KEYINPUT70), .Z(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n437), .A3(new_n436), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT27), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n210), .A2(new_n442), .A3(G210), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n210), .B2(G210), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT26), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n446), .A2(new_n449), .A3(G101), .ZN(new_n450));
  AOI21_X1  g264(.A(G101), .B1(new_n446), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n439), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT31), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n439), .A2(new_n441), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n436), .A2(new_n437), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT73), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT73), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n436), .A2(new_n460), .A3(new_n437), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n440), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n430), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n441), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT28), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n452), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n377), .B1(new_n457), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT74), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(KEYINPUT74), .A3(new_n470), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n469), .B2(new_n470), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n463), .B1(new_n441), .B2(new_n465), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n463), .B2(new_n462), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n454), .B(new_n456), .C1(new_n478), .C2(new_n452), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n377), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n473), .A2(new_n474), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n439), .A2(new_n441), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n452), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT29), .B(new_n484), .C1(new_n452), .C2(new_n478), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n458), .B(new_n440), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT28), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n464), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n452), .A2(KEYINPUT29), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n264), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G472), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n376), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G469), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(new_n264), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n240), .A2(G107), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n240), .A2(G107), .ZN(new_n499));
  OAI21_X1  g313(.A(G101), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT3), .B1(new_n240), .B2(G107), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n302), .A3(G104), .ZN(new_n503));
  INV_X1    g317(.A(G101), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n497), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT1), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n380), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n386), .B2(new_n389), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n387), .A2(G128), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n511), .A2(KEYINPUT10), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n416), .A2(new_n420), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n501), .A2(new_n503), .A3(new_n497), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G101), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT4), .A3(new_n505), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n517), .A3(G101), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n419), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n506), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n433), .A2(KEYINPUT10), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n512), .A2(new_n513), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n513), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n519), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n511), .A2(KEYINPUT10), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n328), .A2(G227), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT80), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT80), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n528), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G110), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n530), .A2(new_n534), .A3(G140), .ZN(new_n535));
  AOI21_X1  g349(.A(G140), .B1(new_n530), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n433), .A2(new_n520), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n523), .B1(new_n540), .B2(new_n511), .ZN(new_n541));
  NOR2_X1   g355(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n523), .B(new_n542), .C1(new_n540), .C2(new_n511), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n522), .A2(new_n545), .A3(new_n537), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n539), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n496), .B1(new_n548), .B2(new_n495), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n522), .A2(new_n545), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n538), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n522), .A2(new_n526), .A3(new_n537), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(G469), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n494), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G224), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT84), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n419), .A2(new_n189), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n400), .A2(new_n189), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n562), .A3(new_n560), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT86), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n516), .A2(new_n430), .A3(new_n518), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT5), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n569), .B(G113), .C1(KEYINPUT5), .C2(new_n424), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n520), .A2(new_n426), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n426), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n506), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n572), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n565), .A2(new_n567), .A3(new_n573), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n561), .A2(new_n562), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n558), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n572), .B1(new_n568), .B2(new_n571), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n573), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT6), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n582), .A2(KEYINPUT83), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT83), .B1(new_n582), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n581), .B(new_n584), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n588), .A3(new_n264), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n579), .A2(new_n588), .A3(new_n264), .A4(new_n590), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G214), .B1(G237), .B2(G902), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n555), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n340), .A2(new_n492), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT33), .B1(new_n316), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n304), .A2(new_n309), .ZN(new_n603));
  INV_X1    g417(.A(new_n313), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n314), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n605), .B(new_n314), .C1(KEYINPUT100), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(G478), .B(new_n264), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n317), .A2(new_n318), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n279), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n594), .A2(new_n595), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n335), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n479), .A2(new_n264), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G472), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n469), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n376), .A2(new_n555), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n269), .B1(new_n268), .B2(new_n264), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n625), .B1(new_n272), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n266), .A2(KEYINPUT101), .A3(new_n270), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n277), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n629), .A2(new_n322), .A3(new_n615), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n357), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n370), .A2(new_n373), .B1(new_n374), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n620), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n340), .A2(new_n598), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT37), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n533), .ZN(G12));
  AOI21_X1  g454(.A(new_n636), .B1(new_n481), .B2(new_n491), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n327), .B1(new_n331), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n629), .A2(new_n322), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n614), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n641), .A2(new_n645), .A3(new_n554), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  XNOR2_X1  g462(.A(new_n643), .B(KEYINPUT39), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n555), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n322), .A3(new_n279), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n264), .B1(new_n486), .B2(new_n452), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n482), .A2(new_n452), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n481), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n636), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n594), .B(KEYINPUT38), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n595), .B(new_n659), .C1(new_n650), .C2(new_n651), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n653), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n205), .ZN(G45));
  AND3_X1   g476(.A1(new_n279), .A2(new_n612), .A3(new_n644), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n641), .A2(new_n663), .A3(new_n554), .A4(new_n646), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  NOR2_X1   g479(.A1(new_n548), .A2(new_n495), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n548), .A2(new_n495), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n493), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n492), .A2(new_n617), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND3_X1  g487(.A1(new_n492), .A2(new_n630), .A3(new_n670), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NAND3_X1  g489(.A1(new_n670), .A2(KEYINPUT102), .A3(new_n646), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n669), .B2(new_n614), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n340), .A2(new_n641), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  AOI21_X1  g495(.A(new_n452), .B1(new_n487), .B2(new_n464), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n377), .B1(new_n682), .B2(new_n457), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n619), .A2(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n375), .A2(new_n684), .A3(new_n615), .A4(new_n670), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n279), .A2(new_n322), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT103), .B1(new_n279), .B2(new_n322), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  INV_X1    g505(.A(new_n636), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n679), .A2(new_n692), .A3(new_n663), .A4(new_n684), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n552), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n551), .A2(new_n552), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n696), .B1(new_n697), .B2(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n494), .B1(new_n699), .B2(new_n549), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n592), .A2(new_n701), .A3(new_n593), .A4(new_n595), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT105), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n663), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n479), .A2(KEYINPUT32), .A3(new_n377), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n491), .A2(new_n471), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n375), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT42), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n492), .A2(new_n711), .A3(new_n663), .A4(new_n705), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n710), .A2(KEYINPUT106), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  NAND3_X1  g532(.A1(new_n492), .A2(new_n645), .A3(new_n705), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  NAND2_X1  g534(.A1(new_n698), .A2(KEYINPUT45), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n697), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(G469), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n496), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n727));
  INV_X1    g541(.A(new_n668), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n727), .B(new_n731), .C1(KEYINPUT46), .C2(new_n726), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n493), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n649), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n704), .A2(new_n702), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n280), .A2(new_n612), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n739), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n620), .B(new_n692), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n734), .B(new_n736), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT109), .B(G137), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G39));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n732), .B2(new_n493), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n481), .A2(new_n376), .A3(new_n491), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n732), .A2(new_n749), .A3(new_n493), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n663), .A2(new_n736), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  NAND3_X1  g571(.A1(new_n736), .A2(KEYINPUT115), .A3(new_n670), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n735), .B2(new_n669), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n327), .C1(new_n740), .C2(new_n742), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n762), .A2(new_n763), .A3(new_n709), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n762), .B2(new_n709), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n376), .B1(new_n758), .B2(new_n760), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n657), .A2(new_n326), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n279), .A3(new_n612), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n323), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n692), .A2(new_n684), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n280), .A3(new_n767), .ZN(new_n771));
  OAI22_X1  g585(.A1(new_n762), .A2(new_n770), .B1(new_n612), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n684), .A2(new_n375), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n670), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n327), .B(new_n774), .C1(new_n740), .C2(new_n742), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT114), .B1(KEYINPUT113), .B2(KEYINPUT50), .ZN(new_n776));
  NOR2_X1   g590(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n659), .A2(new_n595), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n775), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n772), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n740), .A2(new_n742), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n326), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n773), .A3(new_n736), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n728), .A2(new_n666), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n751), .A2(new_n753), .B1(new_n494), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n782), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n769), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(KEYINPUT116), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n494), .ZN(new_n792));
  INV_X1    g606(.A(new_n753), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n750), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(KEYINPUT51), .B(new_n782), .C1(new_n797), .C2(new_n785), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n800));
  INV_X1    g614(.A(new_n322), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n613), .B1(new_n801), .B2(new_n279), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n597), .A2(new_n335), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n621), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n599), .A2(new_n680), .A3(new_n638), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n690), .A2(new_n671), .A3(new_n674), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n627), .A2(new_n628), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n801), .A3(new_n278), .A4(new_n644), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n704), .A2(new_n554), .A3(new_n702), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n481), .B2(new_n491), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n629), .A2(KEYINPUT110), .A3(new_n801), .A4(new_n644), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n663), .A2(new_n705), .A3(new_n684), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n692), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n808), .B1(new_n819), .B2(new_n719), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n636), .B1(new_n816), .B2(new_n817), .ZN(new_n821));
  INV_X1    g635(.A(new_n719), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n821), .A2(KEYINPUT111), .A3(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n717), .B(new_n807), .C1(new_n820), .C2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n647), .A2(new_n664), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n646), .B1(new_n688), .B2(new_n689), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n657), .A2(new_n636), .A3(new_n644), .A4(new_n700), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n825), .A2(new_n828), .A3(KEYINPUT52), .A4(new_n693), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n647), .A2(new_n693), .A3(new_n664), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n826), .A2(new_n827), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n800), .B1(new_n824), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n833), .A2(KEYINPUT112), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n833), .A3(KEYINPUT112), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n805), .A2(new_n713), .A3(new_n806), .A4(new_n800), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n819), .A2(new_n808), .A3(new_n719), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT111), .B1(new_n821), .B2(new_n822), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n784), .A2(new_n679), .A3(new_n773), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT53), .B1(new_n824), .B2(new_n834), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n836), .A2(new_n837), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n848), .B(KEYINPUT54), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n799), .A2(new_n846), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n728), .A2(KEYINPUT49), .A3(new_n666), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT49), .B1(new_n728), .B2(new_n666), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n375), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n657), .A2(new_n659), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n737), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n493), .A3(new_n596), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(G75));
  NOR2_X1   g674(.A1(new_n328), .A2(G952), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT118), .Z(new_n862));
  AOI21_X1  g676(.A(new_n264), .B1(new_n835), .B2(new_n842), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(new_n581), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT117), .B1(new_n843), .B2(G902), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n870), .B(new_n264), .C1(new_n835), .C2(new_n842), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n591), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n868), .B1(new_n872), .B2(new_n874), .ZN(G51));
  NAND2_X1  g689(.A1(new_n539), .A2(new_n547), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n845), .B1(new_n835), .B2(new_n842), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n496), .B(KEYINPUT57), .Z(new_n880));
  OAI21_X1  g694(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n724), .B(KEYINPUT119), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n869), .B2(new_n871), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n861), .B1(new_n881), .B2(new_n883), .ZN(G54));
  AND2_X1   g698(.A1(KEYINPUT58), .A2(G475), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n869), .B2(new_n871), .ZN(new_n886));
  INV_X1    g700(.A(new_n262), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n861), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n262), .B(new_n885), .C1(new_n869), .C2(new_n871), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G60));
  OR2_X1    g705(.A1(new_n606), .A2(new_n609), .ZN(new_n892));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT121), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT120), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT59), .Z(new_n896));
  OAI211_X1 g710(.A(new_n892), .B(new_n896), .C1(new_n877), .C2(new_n878), .ZN(new_n897));
  INV_X1    g711(.A(new_n896), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n846), .B2(new_n851), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n862), .B(new_n897), .C1(new_n899), .C2(new_n892), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(G63));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n371), .B(KEYINPUT60), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n365), .B1(new_n844), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n862), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n635), .B(KEYINPUT122), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n844), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n902), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n908), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n862), .A4(new_n904), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(G66));
  OAI21_X1  g726(.A(G953), .B1(new_n334), .B2(new_n556), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n807), .B2(new_n329), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n865), .B1(G898), .B2(new_n328), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G69));
  NAND2_X1  g730(.A1(new_n422), .A2(new_n438), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n223), .A2(new_n225), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n920));
  NAND2_X1  g734(.A1(G227), .A2(G900), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n329), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n329), .A2(G900), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n735), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n826), .A2(new_n709), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n734), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n756), .A2(new_n693), .A3(new_n825), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n822), .B1(new_n715), .B2(new_n716), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n919), .B(new_n923), .C1(new_n932), .C2(new_n329), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n492), .A2(new_n802), .A3(new_n650), .A4(new_n736), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n831), .A2(new_n661), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n746), .A2(new_n756), .A3(new_n934), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n328), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n919), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n933), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n933), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n922), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n933), .A2(new_n944), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT125), .ZN(new_n950));
  INV_X1    g764(.A(new_n922), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n933), .A2(new_n944), .A3(new_n945), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(new_n953), .ZN(G72));
  XOR2_X1   g768(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n939), .A2(new_n941), .ZN(new_n958));
  INV_X1    g772(.A(new_n807), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n655), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n932), .B2(new_n959), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n482), .A2(new_n452), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n964), .A3(new_n889), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n655), .A3(new_n963), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n967), .B2(new_n957), .ZN(G57));
endmodule


