

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773;

  AND2_X1 U379 ( .A1(n391), .A2(n390), .ZN(n399) );
  AND2_X1 U380 ( .A1(n582), .A2(n654), .ZN(n583) );
  XNOR2_X1 U381 ( .A(n388), .B(n387), .ZN(n771) );
  XNOR2_X1 U382 ( .A(n386), .B(KEYINPUT101), .ZN(n770) );
  INV_X1 U383 ( .A(n562), .ZN(n360) );
  BUF_X1 U384 ( .A(n696), .Z(n358) );
  INV_X1 U385 ( .A(n508), .ZN(n357) );
  XNOR2_X1 U386 ( .A(n521), .B(n367), .ZN(n621) );
  XOR2_X1 U387 ( .A(G143), .B(G128), .Z(n516) );
  NOR2_X2 U388 ( .A1(n613), .A2(n528), .ZN(n530) );
  XNOR2_X2 U389 ( .A(n523), .B(n522), .ZN(n613) );
  XNOR2_X2 U390 ( .A(n506), .B(n505), .ZN(n610) );
  XNOR2_X1 U391 ( .A(n453), .B(n357), .ZN(n363) );
  OR2_X2 U392 ( .A1(n476), .A2(G902), .ZN(n438) );
  INV_X2 U393 ( .A(G953), .ZN(n761) );
  NOR2_X2 U394 ( .A1(n726), .A2(G902), .ZN(n506) );
  INV_X1 U395 ( .A(n510), .ZN(n359) );
  NAND2_X1 U396 ( .A1(n421), .A2(n416), .ZN(n415) );
  AND2_X1 U397 ( .A1(n414), .A2(n366), .ZN(n417) );
  AND2_X1 U398 ( .A1(n413), .A2(n554), .ZN(n416) );
  NOR2_X1 U399 ( .A1(n460), .A2(n401), .ZN(n561) );
  AND2_X1 U400 ( .A1(n579), .A2(n569), .ZN(n567) );
  XNOR2_X1 U401 ( .A(n495), .B(n494), .ZN(n690) );
  XNOR2_X1 U402 ( .A(n432), .B(KEYINPUT3), .ZN(n510) );
  XNOR2_X1 U403 ( .A(G119), .B(G113), .ZN(n432) );
  INV_X1 U404 ( .A(n619), .ZN(n361) );
  BUF_X1 U405 ( .A(n570), .Z(n362) );
  XNOR2_X1 U406 ( .A(n530), .B(n529), .ZN(n570) );
  XNOR2_X1 U407 ( .A(n610), .B(n507), .ZN(n579) );
  BUF_X1 U408 ( .A(n610), .Z(n364) );
  XOR2_X1 U409 ( .A(KEYINPUT70), .B(G131), .Z(n540) );
  XNOR2_X1 U410 ( .A(n482), .B(n405), .ZN(n531) );
  INV_X1 U411 ( .A(KEYINPUT8), .ZN(n405) );
  INV_X1 U412 ( .A(n690), .ZN(n411) );
  XNOR2_X1 U413 ( .A(n553), .B(n552), .ZN(n574) );
  XNOR2_X1 U414 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n541) );
  XOR2_X1 U416 ( .A(G146), .B(G125), .Z(n517) );
  XNOR2_X1 U417 ( .A(G137), .B(G128), .ZN(n480) );
  XNOR2_X1 U418 ( .A(n404), .B(n402), .ZN(n535) );
  XNOR2_X1 U419 ( .A(n549), .B(n758), .ZN(n729) );
  XNOR2_X1 U420 ( .A(n548), .B(n461), .ZN(n549) );
  NOR2_X1 U421 ( .A1(n646), .A2(n647), .ZN(n368) );
  XNOR2_X1 U422 ( .A(KEYINPUT79), .B(KEYINPUT48), .ZN(n644) );
  NAND2_X1 U423 ( .A1(n441), .A2(n444), .ZN(n443) );
  AND2_X1 U424 ( .A1(n448), .A2(KEYINPUT39), .ZN(n444) );
  OR2_X1 U425 ( .A1(n448), .A2(KEYINPUT39), .ZN(n446) );
  XNOR2_X1 U426 ( .A(n558), .B(KEYINPUT22), .ZN(n559) );
  XNOR2_X1 U427 ( .A(n493), .B(n459), .ZN(n494) );
  BUF_X1 U428 ( .A(n726), .Z(n397) );
  NOR2_X1 U429 ( .A1(n641), .A2(KEYINPUT47), .ZN(n394) );
  INV_X1 U430 ( .A(G101), .ZN(n452) );
  XNOR2_X1 U431 ( .A(n465), .B(n359), .ZN(n467) );
  XNOR2_X1 U432 ( .A(n540), .B(G137), .ZN(n462) );
  INV_X1 U433 ( .A(n533), .ZN(n393) );
  NAND2_X1 U434 ( .A1(n531), .A2(G217), .ZN(n404) );
  XNOR2_X1 U435 ( .A(n532), .B(n403), .ZN(n402) );
  INV_X1 U436 ( .A(KEYINPUT95), .ZN(n403) );
  XOR2_X1 U437 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n532) );
  XOR2_X1 U438 ( .A(KEYINPUT93), .B(KEYINPUT12), .Z(n543) );
  XOR2_X1 U439 ( .A(G104), .B(G122), .Z(n547) );
  XNOR2_X1 U440 ( .A(n389), .B(n514), .ZN(n515) );
  XOR2_X1 U441 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n514) );
  XNOR2_X1 U442 ( .A(n513), .B(KEYINPUT17), .ZN(n389) );
  INV_X1 U443 ( .A(n516), .ZN(n518) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n524) );
  NOR2_X1 U445 ( .A1(n434), .A2(n433), .ZN(n645) );
  XNOR2_X1 U446 ( .A(n638), .B(n639), .ZN(n433) );
  NAND2_X1 U447 ( .A1(n629), .A2(n435), .ZN(n434) );
  NOR2_X1 U448 ( .A1(n598), .A2(n449), .ZN(n448) );
  NOR2_X1 U449 ( .A1(G902), .A2(G237), .ZN(n509) );
  XNOR2_X1 U450 ( .A(KEYINPUT85), .B(n475), .ZN(n648) );
  XOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .Z(n475) );
  NOR2_X1 U452 ( .A1(n570), .A2(n425), .ZN(n420) );
  XOR2_X1 U453 ( .A(G107), .B(G104), .Z(n496) );
  XNOR2_X1 U454 ( .A(n632), .B(KEYINPUT107), .ZN(n633) );
  NAND2_X1 U455 ( .A1(n362), .A2(n425), .ZN(n423) );
  INV_X1 U456 ( .A(KEYINPUT100), .ZN(n409) );
  INV_X1 U457 ( .A(KEYINPUT32), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n609), .B(n395), .ZN(n611) );
  XNOR2_X1 U459 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n395) );
  INV_X1 U460 ( .A(G472), .ZN(n437) );
  XNOR2_X1 U461 ( .A(n489), .B(n758), .ZN(n736) );
  NAND2_X1 U462 ( .A1(n368), .A2(n746), .ZN(n678) );
  NAND2_X1 U463 ( .A1(n442), .A2(n443), .ZN(n630) );
  INV_X1 U464 ( .A(n445), .ZN(n442) );
  NOR2_X1 U465 ( .A1(n440), .A2(n445), .ZN(n631) );
  NAND2_X1 U466 ( .A1(n443), .A2(n663), .ZN(n440) );
  AND2_X1 U467 ( .A1(n563), .A2(n455), .ZN(n454) );
  INV_X1 U468 ( .A(KEYINPUT122), .ZN(n378) );
  INV_X1 U469 ( .A(KEYINPUT60), .ZN(n380) );
  XNOR2_X1 U470 ( .A(n397), .B(n725), .ZN(n400) );
  AND2_X1 U471 ( .A1(n563), .A2(n408), .ZN(n365) );
  OR2_X1 U472 ( .A1(n616), .A2(KEYINPUT35), .ZN(n366) );
  AND2_X1 U473 ( .A1(n520), .A2(G210), .ZN(n367) );
  AND2_X1 U474 ( .A1(n420), .A2(n419), .ZN(n369) );
  INV_X1 U475 ( .A(KEYINPUT39), .ZN(n450) );
  XOR2_X1 U476 ( .A(n476), .B(KEYINPUT62), .Z(n370) );
  XOR2_X1 U477 ( .A(n732), .B(n731), .Z(n371) );
  XOR2_X1 U478 ( .A(n729), .B(n728), .Z(n372) );
  OR2_X1 U479 ( .A1(n650), .A2(n648), .ZN(n373) );
  XOR2_X1 U480 ( .A(n722), .B(n721), .Z(n374) );
  NOR2_X1 U481 ( .A1(G952), .A2(n761), .ZN(n740) );
  INV_X1 U482 ( .A(n740), .ZN(n390) );
  XNOR2_X1 U483 ( .A(n724), .B(n400), .ZN(n727) );
  AND2_X2 U484 ( .A1(n430), .A2(n428), .ZN(n375) );
  AND2_X1 U485 ( .A1(n430), .A2(n428), .ZN(n734) );
  NAND2_X1 U486 ( .A1(n500), .A2(n451), .ZN(n406) );
  XNOR2_X1 U487 ( .A(n412), .B(n759), .ZN(n726) );
  XNOR2_X1 U488 ( .A(n406), .B(n503), .ZN(n412) );
  XNOR2_X1 U489 ( .A(n376), .B(n377), .ZN(G57) );
  NAND2_X1 U490 ( .A1(n396), .A2(n390), .ZN(n376) );
  XOR2_X1 U491 ( .A(n653), .B(n652), .Z(n377) );
  XNOR2_X1 U492 ( .A(n379), .B(n378), .ZN(G63) );
  NAND2_X1 U493 ( .A1(n384), .A2(n390), .ZN(n379) );
  XNOR2_X1 U494 ( .A(n381), .B(n380), .ZN(G60) );
  NAND2_X1 U495 ( .A1(n385), .A2(n390), .ZN(n381) );
  BUF_X1 U496 ( .A(n579), .Z(n401) );
  INV_X1 U497 ( .A(n401), .ZN(n455) );
  NOR2_X1 U498 ( .A1(n771), .A2(n770), .ZN(n382) );
  NOR2_X1 U499 ( .A1(n771), .A2(n770), .ZN(n407) );
  XNOR2_X1 U500 ( .A(n383), .B(KEYINPUT44), .ZN(n586) );
  NAND2_X1 U501 ( .A1(n564), .A2(n407), .ZN(n383) );
  XNOR2_X1 U502 ( .A(n733), .B(n371), .ZN(n384) );
  XNOR2_X1 U503 ( .A(n730), .B(n372), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n360), .A2(n561), .ZN(n386) );
  NAND2_X1 U505 ( .A1(n431), .A2(n373), .ZN(n430) );
  AND2_X2 U506 ( .A1(n418), .A2(n417), .ZN(n398) );
  INV_X1 U507 ( .A(KEYINPUT67), .ZN(n470) );
  NOR2_X1 U508 ( .A1(n649), .A2(n648), .ZN(n588) );
  XNOR2_X1 U509 ( .A(n587), .B(KEYINPUT45), .ZN(n649) );
  NAND2_X1 U510 ( .A1(n360), .A2(n365), .ZN(n388) );
  NAND2_X2 U511 ( .A1(n398), .A2(n415), .ZN(n565) );
  XNOR2_X1 U512 ( .A(n723), .B(n374), .ZN(n391) );
  NAND2_X1 U513 ( .A1(n511), .A2(n392), .ZN(n512) );
  NAND2_X1 U514 ( .A1(n359), .A2(n393), .ZN(n392) );
  NOR2_X1 U515 ( .A1(n394), .A2(KEYINPUT77), .ZN(n642) );
  XNOR2_X1 U516 ( .A(n537), .B(n462), .ZN(n504) );
  NOR2_X1 U517 ( .A1(n643), .A2(n436), .ZN(n435) );
  INV_X1 U518 ( .A(n746), .ZN(n426) );
  XNOR2_X1 U519 ( .A(n651), .B(n370), .ZN(n396) );
  XNOR2_X1 U520 ( .A(n458), .B(n519), .ZN(n457) );
  NAND2_X1 U521 ( .A1(n621), .A2(n679), .ZN(n523) );
  XNOR2_X1 U522 ( .A(n741), .B(n457), .ZN(n456) );
  XNOR2_X1 U523 ( .A(n399), .B(KEYINPUT56), .ZN(G51) );
  AND2_X2 U524 ( .A1(n565), .A2(KEYINPUT68), .ZN(n564) );
  XNOR2_X1 U525 ( .A(n406), .B(n456), .ZN(n720) );
  NAND2_X1 U526 ( .A1(n566), .A2(n382), .ZN(n584) );
  XNOR2_X1 U527 ( .A(n410), .B(n409), .ZN(n408) );
  NAND2_X1 U528 ( .A1(n401), .A2(n411), .ZN(n410) );
  NAND2_X1 U529 ( .A1(n363), .A2(n369), .ZN(n414) );
  NAND2_X1 U530 ( .A1(n363), .A2(n420), .ZN(n413) );
  NAND2_X1 U531 ( .A1(n422), .A2(n419), .ZN(n418) );
  AND2_X1 U532 ( .A1(n616), .A2(KEYINPUT35), .ZN(n419) );
  INV_X1 U533 ( .A(n422), .ZN(n421) );
  NAND2_X1 U534 ( .A1(n424), .A2(n423), .ZN(n422) );
  NAND2_X1 U535 ( .A1(n713), .A2(n425), .ZN(n424) );
  INV_X1 U536 ( .A(KEYINPUT34), .ZN(n425) );
  NOR2_X1 U537 ( .A1(n426), .A2(n650), .ZN(n429) );
  NAND2_X1 U538 ( .A1(n427), .A2(n368), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n588), .B(KEYINPUT78), .ZN(n427) );
  NAND2_X1 U540 ( .A1(n368), .A2(n429), .ZN(n428) );
  NAND2_X1 U541 ( .A1(n640), .A2(n773), .ZN(n436) );
  XNOR2_X2 U542 ( .A(n438), .B(n437), .ZN(n571) );
  XNOR2_X1 U543 ( .A(n439), .B(n468), .ZN(n476) );
  XNOR2_X1 U544 ( .A(n504), .B(n498), .ZN(n439) );
  INV_X1 U545 ( .A(n597), .ZN(n441) );
  NAND2_X1 U546 ( .A1(n447), .A2(n446), .ZN(n445) );
  NAND2_X1 U547 ( .A1(n597), .A2(n450), .ZN(n447) );
  NOR2_X1 U548 ( .A1(n597), .A2(n598), .ZN(n617) );
  INV_X1 U549 ( .A(n680), .ZN(n449) );
  INV_X1 U550 ( .A(n498), .ZN(n499) );
  NAND2_X1 U551 ( .A1(n498), .A2(n497), .ZN(n451) );
  XNOR2_X2 U552 ( .A(n474), .B(n452), .ZN(n498) );
  XNOR2_X2 U553 ( .A(n453), .B(n508), .ZN(n713) );
  NAND2_X1 U554 ( .A1(n567), .A2(n602), .ZN(n453) );
  NAND2_X1 U555 ( .A1(n360), .A2(n454), .ZN(n580) );
  INV_X1 U556 ( .A(n515), .ZN(n458) );
  XNOR2_X2 U557 ( .A(n512), .B(KEYINPUT16), .ZN(n741) );
  XOR2_X1 U558 ( .A(n492), .B(n491), .Z(n459) );
  OR2_X1 U559 ( .A1(n358), .A2(n690), .ZN(n460) );
  XOR2_X1 U560 ( .A(n547), .B(n546), .Z(n461) );
  INV_X1 U561 ( .A(G475), .ZN(n550) );
  INV_X1 U562 ( .A(G140), .ZN(n487) );
  INV_X1 U563 ( .A(KEYINPUT41), .ZN(n632) );
  XNOR2_X1 U564 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n507) );
  XNOR2_X1 U565 ( .A(n488), .B(n487), .ZN(n758) );
  XNOR2_X1 U566 ( .A(n599), .B(n361), .ZN(n680) );
  INV_X1 U567 ( .A(KEYINPUT19), .ZN(n522) );
  XNOR2_X1 U568 ( .A(n634), .B(n633), .ZN(n712) );
  XOR2_X1 U569 ( .A(n575), .B(KEYINPUT97), .Z(n667) );
  XOR2_X1 U570 ( .A(G134), .B(n516), .Z(n537) );
  XOR2_X1 U571 ( .A(G116), .B(KEYINPUT5), .Z(n464) );
  XNOR2_X1 U572 ( .A(G146), .B(KEYINPUT74), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U574 ( .A1(n541), .A2(G210), .ZN(n466) );
  XNOR2_X1 U575 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X2 U576 ( .A(KEYINPUT4), .B(KEYINPUT69), .ZN(n469) );
  XNOR2_X2 U577 ( .A(n469), .B(KEYINPUT64), .ZN(n757) );
  INV_X1 U578 ( .A(n757), .ZN(n471) );
  NAND2_X1 U579 ( .A1(n471), .A2(n470), .ZN(n473) );
  NAND2_X1 U580 ( .A1(n757), .A2(KEYINPUT67), .ZN(n472) );
  NAND2_X1 U581 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U582 ( .A(KEYINPUT102), .B(KEYINPUT33), .Z(n508) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(KEYINPUT98), .ZN(n477) );
  INV_X2 U584 ( .A(n571), .ZN(n696) );
  XOR2_X1 U585 ( .A(n477), .B(n696), .Z(n602) );
  NAND2_X1 U586 ( .A1(n648), .A2(G234), .ZN(n478) );
  XNOR2_X1 U587 ( .A(n478), .B(KEYINPUT20), .ZN(n490) );
  NAND2_X1 U588 ( .A1(n490), .A2(G221), .ZN(n479) );
  XOR2_X1 U589 ( .A(n479), .B(KEYINPUT21), .Z(n691) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n481) );
  XNOR2_X1 U591 ( .A(n481), .B(n480), .ZN(n486) );
  XOR2_X1 U592 ( .A(G119), .B(G110), .Z(n484) );
  NAND2_X1 U593 ( .A1(G234), .A2(n761), .ZN(n482) );
  NAND2_X1 U594 ( .A1(G221), .A2(n531), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n489) );
  XNOR2_X1 U597 ( .A(n517), .B(KEYINPUT10), .ZN(n488) );
  NOR2_X1 U598 ( .A1(G902), .A2(n736), .ZN(n495) );
  NAND2_X1 U599 ( .A1(n490), .A2(G217), .ZN(n493) );
  XOR2_X1 U600 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n492) );
  XNOR2_X1 U601 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n491) );
  NAND2_X1 U602 ( .A1(n691), .A2(n690), .ZN(n698) );
  INV_X1 U603 ( .A(n698), .ZN(n569) );
  XNOR2_X1 U604 ( .A(G110), .B(n496), .ZN(n743) );
  INV_X1 U605 ( .A(n743), .ZN(n497) );
  NAND2_X1 U606 ( .A1(n499), .A2(n743), .ZN(n500) );
  XOR2_X1 U607 ( .A(G146), .B(G140), .Z(n502) );
  NAND2_X1 U608 ( .A1(G227), .A2(n761), .ZN(n501) );
  XNOR2_X1 U609 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U610 ( .A(n504), .B(KEYINPUT88), .ZN(n759) );
  XNOR2_X1 U611 ( .A(KEYINPUT71), .B(G469), .ZN(n505) );
  XNOR2_X1 U612 ( .A(n509), .B(KEYINPUT73), .ZN(n520) );
  NAND2_X1 U613 ( .A1(G214), .A2(n520), .ZN(n679) );
  XOR2_X1 U614 ( .A(G116), .B(G122), .Z(n533) );
  NAND2_X1 U615 ( .A1(n510), .A2(n533), .ZN(n511) );
  NAND2_X1 U616 ( .A1(G224), .A2(n761), .ZN(n513) );
  XOR2_X1 U617 ( .A(n518), .B(n517), .Z(n519) );
  NAND2_X1 U618 ( .A1(n720), .A2(n648), .ZN(n521) );
  XNOR2_X1 U619 ( .A(n524), .B(KEYINPUT14), .ZN(n525) );
  NAND2_X1 U620 ( .A1(G952), .A2(n525), .ZN(n711) );
  NOR2_X1 U621 ( .A1(G953), .A2(n711), .ZN(n593) );
  NAND2_X1 U622 ( .A1(G902), .A2(n525), .ZN(n589) );
  XOR2_X1 U623 ( .A(G898), .B(KEYINPUT86), .Z(n751) );
  NAND2_X1 U624 ( .A1(G953), .A2(n751), .ZN(n745) );
  NOR2_X1 U625 ( .A1(n589), .A2(n745), .ZN(n526) );
  XOR2_X1 U626 ( .A(KEYINPUT87), .B(n526), .Z(n527) );
  NOR2_X1 U627 ( .A1(n593), .A2(n527), .ZN(n528) );
  XNOR2_X1 U628 ( .A(KEYINPUT83), .B(KEYINPUT0), .ZN(n529) );
  XNOR2_X1 U629 ( .A(G107), .B(n533), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U631 ( .A(n537), .B(n536), .ZN(n732) );
  NOR2_X1 U632 ( .A1(G902), .A2(n732), .ZN(n539) );
  XNOR2_X1 U633 ( .A(KEYINPUT96), .B(G478), .ZN(n538) );
  XNOR2_X1 U634 ( .A(n539), .B(n538), .ZN(n577) );
  XNOR2_X1 U635 ( .A(n540), .B(KEYINPUT11), .ZN(n545) );
  NAND2_X1 U636 ( .A1(G214), .A2(n541), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U638 ( .A(n545), .B(n544), .ZN(n548) );
  XNOR2_X1 U639 ( .A(G143), .B(G113), .ZN(n546) );
  NOR2_X1 U640 ( .A1(G902), .A2(n729), .ZN(n553) );
  XNOR2_X1 U641 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n551) );
  NOR2_X1 U642 ( .A1(n577), .A2(n574), .ZN(n616) );
  INV_X1 U643 ( .A(KEYINPUT35), .ZN(n554) );
  INV_X1 U644 ( .A(n691), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n577), .A2(n574), .ZN(n682) );
  NOR2_X1 U646 ( .A1(n555), .A2(n682), .ZN(n556) );
  XNOR2_X1 U647 ( .A(n556), .B(KEYINPUT99), .ZN(n557) );
  NOR2_X1 U648 ( .A1(n570), .A2(n557), .ZN(n560) );
  XNOR2_X1 U649 ( .A(KEYINPUT65), .B(KEYINPUT72), .ZN(n558) );
  XNOR2_X1 U650 ( .A(n560), .B(n559), .ZN(n562) );
  INV_X1 U651 ( .A(n602), .ZN(n563) );
  NOR2_X1 U652 ( .A1(KEYINPUT68), .A2(n565), .ZN(n566) );
  NAND2_X1 U653 ( .A1(n358), .A2(n567), .ZN(n703) );
  NOR2_X1 U654 ( .A1(n703), .A2(n362), .ZN(n568) );
  XNOR2_X1 U655 ( .A(n568), .B(KEYINPUT31), .ZN(n669) );
  NAND2_X1 U656 ( .A1(n364), .A2(n569), .ZN(n598) );
  NOR2_X1 U657 ( .A1(n362), .A2(n598), .ZN(n572) );
  NAND2_X1 U658 ( .A1(n572), .A2(n571), .ZN(n656) );
  NAND2_X1 U659 ( .A1(n669), .A2(n656), .ZN(n573) );
  XNOR2_X1 U660 ( .A(n573), .B(KEYINPUT92), .ZN(n578) );
  INV_X1 U661 ( .A(n574), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n576), .A2(n577), .ZN(n575) );
  NOR2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n660) );
  INV_X1 U664 ( .A(n660), .ZN(n670) );
  NAND2_X1 U665 ( .A1(n667), .A2(n670), .ZN(n607) );
  NAND2_X1 U666 ( .A1(n578), .A2(n607), .ZN(n582) );
  XNOR2_X1 U667 ( .A(KEYINPUT81), .B(n580), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n581), .A2(n690), .ZN(n654) );
  NAND2_X1 U669 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n587) );
  OR2_X1 U671 ( .A1(n761), .A2(n589), .ZN(n590) );
  XOR2_X1 U672 ( .A(KEYINPUT103), .B(n590), .Z(n591) );
  NOR2_X1 U673 ( .A1(G900), .A2(n591), .ZN(n592) );
  NOR2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U675 ( .A(KEYINPUT76), .B(n594), .Z(n600) );
  NAND2_X1 U676 ( .A1(n696), .A2(n679), .ZN(n595) );
  XOR2_X1 U677 ( .A(KEYINPUT30), .B(n595), .Z(n596) );
  NAND2_X1 U678 ( .A1(n600), .A2(n596), .ZN(n597) );
  INV_X1 U679 ( .A(KEYINPUT38), .ZN(n599) );
  OR2_X1 U680 ( .A1(n670), .A2(n630), .ZN(n676) );
  INV_X1 U681 ( .A(n667), .ZN(n663) );
  NAND2_X1 U682 ( .A1(n600), .A2(n691), .ZN(n601) );
  NOR2_X1 U683 ( .A1(n690), .A2(n601), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n663), .A2(n608), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n679), .A2(n602), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n622) );
  NAND2_X1 U687 ( .A1(n622), .A2(n455), .ZN(n605) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT43), .ZN(n606) );
  INV_X1 U689 ( .A(n621), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n606), .A2(n619), .ZN(n677) );
  NAND2_X1 U691 ( .A1(n676), .A2(n677), .ZN(n647) );
  INV_X1 U692 ( .A(n607), .ZN(n684) );
  INV_X1 U693 ( .A(KEYINPUT77), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n684), .A2(n626), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n608), .A2(n696), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n611), .A2(n364), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n612), .B(KEYINPUT106), .ZN(n635) );
  NOR2_X1 U698 ( .A1(n635), .A2(n613), .ZN(n664) );
  NAND2_X1 U699 ( .A1(n614), .A2(n664), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n615), .A2(KEYINPUT47), .ZN(n640) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U703 ( .A(KEYINPUT104), .B(n620), .Z(n773) );
  XOR2_X1 U704 ( .A(KEYINPUT36), .B(KEYINPUT109), .Z(n624) );
  NAND2_X1 U705 ( .A1(n622), .A2(n361), .ZN(n623) );
  XNOR2_X1 U706 ( .A(n624), .B(n623), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n625), .A2(n455), .ZN(n673) );
  XNOR2_X1 U708 ( .A(n673), .B(KEYINPUT80), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n626), .A2(KEYINPUT47), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  INV_X1 U711 ( .A(KEYINPUT46), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT40), .ZN(n772) );
  XNOR2_X1 U713 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n680), .A2(n679), .ZN(n685) );
  NOR2_X1 U715 ( .A1(n682), .A2(n685), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n712), .A2(n635), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n637), .B(n636), .ZN(n769) );
  NOR2_X1 U718 ( .A1(n772), .A2(n769), .ZN(n638) );
  INV_X1 U719 ( .A(n664), .ZN(n641) );
  NOR2_X1 U720 ( .A1(n684), .A2(n642), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(n646) );
  INV_X1 U722 ( .A(KEYINPUT2), .ZN(n650) );
  INV_X1 U723 ( .A(n649), .ZN(n746) );
  NAND2_X1 U724 ( .A1(n375), .A2(G472), .ZN(n651) );
  XOR2_X1 U725 ( .A(KEYINPUT82), .B(KEYINPUT110), .Z(n653) );
  XNOR2_X1 U726 ( .A(KEYINPUT84), .B(KEYINPUT63), .ZN(n652) );
  XNOR2_X1 U727 ( .A(G101), .B(n654), .ZN(G3) );
  NOR2_X1 U728 ( .A1(n667), .A2(n656), .ZN(n655) );
  XOR2_X1 U729 ( .A(G104), .B(n655), .Z(G6) );
  NOR2_X1 U730 ( .A1(n670), .A2(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(G107), .B(n659), .ZN(G9) );
  XOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  NAND2_X1 U735 ( .A1(n664), .A2(n660), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(G30) );
  XOR2_X1 U737 ( .A(G146), .B(KEYINPUT111), .Z(n666) );
  NAND2_X1 U738 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(G48) );
  NOR2_X1 U740 ( .A1(n667), .A2(n669), .ZN(n668) );
  XOR2_X1 U741 ( .A(G113), .B(n668), .Z(G15) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT112), .B(n671), .Z(n672) );
  XNOR2_X1 U744 ( .A(G116), .B(n672), .ZN(G18) );
  XNOR2_X1 U745 ( .A(G125), .B(n673), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U747 ( .A(G134), .B(KEYINPUT113), .Z(n675) );
  XNOR2_X1 U748 ( .A(n676), .B(n675), .ZN(G36) );
  XNOR2_X1 U749 ( .A(G140), .B(n677), .ZN(G42) );
  XOR2_X1 U750 ( .A(KEYINPUT2), .B(n678), .Z(n717) );
  NOR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n683), .B(KEYINPUT118), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U756 ( .A(KEYINPUT119), .B(n688), .Z(n689) );
  NOR2_X1 U757 ( .A1(n713), .A2(n689), .ZN(n708) );
  XOR2_X1 U758 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n693) );
  OR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n694), .B(KEYINPUT114), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n358), .A2(n695), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT116), .ZN(n702) );
  XOR2_X1 U764 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n700) );
  NAND2_X1 U765 ( .A1(n455), .A2(n698), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U769 ( .A(KEYINPUT51), .B(n705), .ZN(n706) );
  NOR2_X1 U770 ( .A1(n712), .A2(n706), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n709), .B(KEYINPUT52), .ZN(n710) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U775 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U776 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U777 ( .A1(n718), .A2(G953), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n719), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U779 ( .A1(n734), .A2(G210), .ZN(n723) );
  INV_X1 U780 ( .A(n720), .ZN(n722) );
  XOR2_X1 U781 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n721) );
  XOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n725) );
  NAND2_X1 U783 ( .A1(n375), .A2(G469), .ZN(n724) );
  NOR2_X1 U784 ( .A1(n740), .A2(n727), .ZN(G54) );
  NAND2_X1 U785 ( .A1(n375), .A2(G475), .ZN(n730) );
  XOR2_X1 U786 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n728) );
  NAND2_X1 U787 ( .A1(n375), .A2(G478), .ZN(n733) );
  INV_X1 U788 ( .A(KEYINPUT121), .ZN(n731) );
  NAND2_X1 U789 ( .A1(n375), .A2(G217), .ZN(n738) );
  INV_X1 U790 ( .A(KEYINPUT123), .ZN(n735) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(G66) );
  XOR2_X1 U794 ( .A(n741), .B(G101), .Z(n742) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(n744) );
  NAND2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n755) );
  NAND2_X1 U797 ( .A1(n746), .A2(n761), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n747), .B(KEYINPUT125), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n749) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U804 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U805 ( .A(KEYINPUT126), .B(n756), .ZN(G69) );
  XOR2_X1 U806 ( .A(n758), .B(n757), .Z(n760) );
  XNOR2_X1 U807 ( .A(n760), .B(n759), .ZN(n763) );
  XOR2_X1 U808 ( .A(n368), .B(n763), .Z(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n768) );
  XNOR2_X1 U810 ( .A(G227), .B(n763), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U812 ( .A1(G953), .A2(n765), .ZN(n766) );
  XOR2_X1 U813 ( .A(KEYINPUT127), .B(n766), .Z(n767) );
  NAND2_X1 U814 ( .A1(n768), .A2(n767), .ZN(G72) );
  XNOR2_X1 U815 ( .A(n565), .B(G122), .ZN(G24) );
  XOR2_X1 U816 ( .A(G137), .B(n769), .Z(G39) );
  XOR2_X1 U817 ( .A(n770), .B(G110), .Z(G12) );
  XOR2_X1 U818 ( .A(n771), .B(G119), .Z(G21) );
  XOR2_X1 U819 ( .A(n772), .B(G131), .Z(G33) );
  XNOR2_X1 U820 ( .A(G143), .B(n773), .ZN(G45) );
endmodule

