

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(KEYINPUT31), .ZN(n652) );
  AND2_X1 U553 ( .A1(n595), .A2(n686), .ZN(n596) );
  AND2_X1 U554 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U555 ( .A1(n656), .A2(G8), .ZN(n745) );
  INV_X1 U556 ( .A(KEYINPUT99), .ZN(n682) );
  AND2_X1 U557 ( .A1(n521), .A2(G2104), .ZN(n881) );
  NOR2_X1 U558 ( .A1(n554), .A2(G651), .ZN(n791) );
  NOR2_X1 U559 ( .A1(n526), .A2(n525), .ZN(G160) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n517), .Z(n882) );
  NAND2_X1 U562 ( .A1(n882), .A2(G137), .ZN(n520) );
  INV_X1 U563 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U564 ( .A1(G101), .A2(n881), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U566 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n521), .ZN(n877) );
  NAND2_X1 U568 ( .A1(n877), .A2(G125), .ZN(n524) );
  NAND2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U570 ( .A(n522), .B(KEYINPUT68), .Z(n878) );
  NAND2_X1 U571 ( .A1(G113), .A2(n878), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n554) );
  INV_X1 U574 ( .A(G651), .ZN(n534) );
  NOR2_X1 U575 ( .A1(n554), .A2(n534), .ZN(n784) );
  NAND2_X1 U576 ( .A1(G76), .A2(n784), .ZN(n531) );
  XOR2_X1 U577 ( .A(KEYINPUT75), .B(KEYINPUT4), .Z(n529) );
  NOR2_X1 U578 ( .A1(G543), .A2(G651), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT67), .B(n527), .Z(n787) );
  NAND2_X1 U580 ( .A1(G89), .A2(n787), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U583 ( .A(n532), .B(KEYINPUT5), .ZN(n533) );
  XNOR2_X1 U584 ( .A(KEYINPUT76), .B(n533), .ZN(n541) );
  XNOR2_X1 U585 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n539) );
  NAND2_X1 U586 ( .A1(G51), .A2(n791), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n535), .Z(n783) );
  NAND2_X1 U589 ( .A1(G63), .A2(n783), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U593 ( .A(n542), .B(KEYINPUT7), .ZN(n543) );
  XNOR2_X1 U594 ( .A(KEYINPUT78), .B(n543), .ZN(G168) );
  XOR2_X1 U595 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U596 ( .A1(n881), .A2(G102), .ZN(n544) );
  XNOR2_X1 U597 ( .A(n544), .B(KEYINPUT86), .ZN(n546) );
  NAND2_X1 U598 ( .A1(G138), .A2(n882), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n877), .A2(G126), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G114), .A2(n878), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n550), .A2(n549), .ZN(G164) );
  NAND2_X1 U604 ( .A1(G49), .A2(n791), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G74), .A2(G651), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U607 ( .A1(n783), .A2(n553), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n554), .A2(G87), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n556), .A2(n555), .ZN(G288) );
  NAND2_X1 U610 ( .A1(G64), .A2(n783), .ZN(n557) );
  XOR2_X1 U611 ( .A(KEYINPUT70), .B(n557), .Z(n564) );
  NAND2_X1 U612 ( .A1(G90), .A2(n787), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G77), .A2(n784), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G52), .A2(n791), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U618 ( .A1(n564), .A2(n563), .ZN(G171) );
  NAND2_X1 U619 ( .A1(G91), .A2(n787), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G78), .A2(n784), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U622 ( .A1(n783), .A2(G65), .ZN(n567) );
  XOR2_X1 U623 ( .A(KEYINPUT72), .B(n567), .Z(n568) );
  NOR2_X1 U624 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n791), .A2(G53), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n571), .A2(n570), .ZN(G299) );
  NAND2_X1 U627 ( .A1(G88), .A2(n787), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT84), .ZN(n579) );
  NAND2_X1 U629 ( .A1(G50), .A2(n791), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G75), .A2(n784), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U632 ( .A1(G62), .A2(n783), .ZN(n575) );
  XNOR2_X1 U633 ( .A(KEYINPUT83), .B(n575), .ZN(n576) );
  NOR2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G61), .A2(n783), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G86), .A2(n787), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U639 ( .A(KEYINPUT82), .B(n582), .ZN(n585) );
  NAND2_X1 U640 ( .A1(n784), .A2(G73), .ZN(n583) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n583), .Z(n584) );
  NOR2_X1 U642 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n791), .A2(G48), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G85), .A2(n787), .ZN(n589) );
  NAND2_X1 U646 ( .A1(G72), .A2(n784), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U648 ( .A1(G47), .A2(n791), .ZN(n590) );
  XNOR2_X1 U649 ( .A(KEYINPUT69), .B(n590), .ZN(n591) );
  NOR2_X1 U650 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U651 ( .A1(n783), .A2(G60), .ZN(n593) );
  NAND2_X1 U652 ( .A1(n594), .A2(n593), .ZN(G290) );
  INV_X1 U653 ( .A(G303), .ZN(G166) );
  AND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n595) );
  NOR2_X1 U655 ( .A1(G164), .A2(G1384), .ZN(n686) );
  XNOR2_X2 U656 ( .A(n596), .B(KEYINPUT64), .ZN(n629) );
  INV_X1 U657 ( .A(n629), .ZN(n656) );
  NOR2_X1 U658 ( .A1(G1976), .A2(G288), .ZN(n674) );
  NAND2_X1 U659 ( .A1(n674), .A2(KEYINPUT33), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n745), .A2(n597), .ZN(n681) );
  XNOR2_X1 U661 ( .A(G2078), .B(KEYINPUT25), .ZN(n971) );
  NAND2_X1 U662 ( .A1(n629), .A2(n971), .ZN(n599) );
  INV_X1 U663 ( .A(G1961), .ZN(n850) );
  NAND2_X1 U664 ( .A1(n656), .A2(n850), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n649) );
  NAND2_X1 U666 ( .A1(n649), .A2(G171), .ZN(n645) );
  XNOR2_X1 U667 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n643) );
  INV_X1 U668 ( .A(G299), .ZN(n799) );
  NAND2_X1 U669 ( .A1(G2072), .A2(n629), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT27), .ZN(n602) );
  INV_X1 U671 ( .A(G1956), .ZN(n941) );
  NOR2_X1 U672 ( .A1(n629), .A2(n941), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n799), .A2(n604), .ZN(n603) );
  XOR2_X1 U675 ( .A(n603), .B(KEYINPUT28), .Z(n641) );
  NAND2_X1 U676 ( .A1(n799), .A2(n604), .ZN(n639) );
  NAND2_X1 U677 ( .A1(G1996), .A2(n629), .ZN(n606) );
  XNOR2_X1 U678 ( .A(KEYINPUT66), .B(KEYINPUT26), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n606), .B(n605), .ZN(n619) );
  NAND2_X1 U680 ( .A1(G56), .A2(n783), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n607), .Z(n613) );
  NAND2_X1 U682 ( .A1(n787), .A2(G81), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G68), .A2(n784), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT13), .B(n611), .Z(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n791), .A2(G43), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n934) );
  INV_X1 U690 ( .A(G1341), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n629), .A2(n616), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n934), .A2(n617), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n635) );
  NAND2_X1 U694 ( .A1(G66), .A2(n783), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G92), .A2(n787), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G54), .A2(n791), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G79), .A2(n784), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT73), .B(n624), .Z(n625) );
  NOR2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(KEYINPUT15), .B(n627), .ZN(n920) );
  NOR2_X1 U703 ( .A1(n635), .A2(n920), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT95), .ZN(n634) );
  NAND2_X1 U705 ( .A1(G2067), .A2(n629), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n656), .A2(G1348), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U708 ( .A(KEYINPUT96), .B(n632), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n635), .A2(n920), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n655) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n745), .ZN(n668) );
  NOR2_X1 U717 ( .A1(n656), .A2(G2084), .ZN(n665) );
  NOR2_X1 U718 ( .A1(n668), .A2(n665), .ZN(n646) );
  NAND2_X1 U719 ( .A1(G8), .A2(n646), .ZN(n647) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n647), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n648), .A2(G168), .ZN(n651) );
  NOR2_X1 U722 ( .A1(G171), .A2(n649), .ZN(n650) );
  NOR2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n666) );
  NAND2_X1 U726 ( .A1(n666), .A2(G286), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n656), .A2(G2090), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT98), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n745), .A2(G1971), .ZN(n658) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n660), .A2(G303), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U733 ( .A1(G8), .A2(n663), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT32), .ZN(n672) );
  NAND2_X1 U735 ( .A1(G8), .A2(n665), .ZN(n670) );
  INV_X1 U736 ( .A(n666), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n743) );
  NOR2_X1 U740 ( .A1(G1971), .A2(G303), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n918) );
  NAND2_X1 U742 ( .A1(n743), .A2(n918), .ZN(n677) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n915) );
  INV_X1 U744 ( .A(n915), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n745), .A2(n675), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT65), .B(n678), .Z(n679) );
  NOR2_X1 U747 ( .A1(KEYINPUT33), .A2(n679), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n724) );
  XOR2_X1 U750 ( .A(G1981), .B(KEYINPUT100), .Z(n684) );
  XNOR2_X1 U751 ( .A(G305), .B(n684), .ZN(n928) );
  NAND2_X1 U752 ( .A1(G160), .A2(G40), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n736) );
  XNOR2_X1 U754 ( .A(KEYINPUT37), .B(G2067), .ZN(n725) );
  NAND2_X1 U755 ( .A1(n881), .A2(G104), .ZN(n687) );
  XNOR2_X1 U756 ( .A(KEYINPUT87), .B(n687), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n882), .A2(G140), .ZN(n688) );
  XOR2_X1 U758 ( .A(n688), .B(KEYINPUT88), .Z(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U760 ( .A(KEYINPUT89), .B(n691), .Z(n692) );
  XNOR2_X1 U761 ( .A(KEYINPUT34), .B(n692), .ZN(n698) );
  XNOR2_X1 U762 ( .A(KEYINPUT35), .B(KEYINPUT90), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n877), .A2(G128), .ZN(n694) );
  NAND2_X1 U764 ( .A1(G116), .A2(n878), .ZN(n693) );
  NAND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U768 ( .A(n699), .B(KEYINPUT36), .Z(n867) );
  NOR2_X1 U769 ( .A1(n725), .A2(n867), .ZN(n998) );
  NAND2_X1 U770 ( .A1(n736), .A2(n998), .ZN(n733) );
  NAND2_X1 U771 ( .A1(G105), .A2(n881), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n700), .B(KEYINPUT38), .ZN(n708) );
  NAND2_X1 U773 ( .A1(G129), .A2(n877), .ZN(n701) );
  XNOR2_X1 U774 ( .A(n701), .B(KEYINPUT92), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n882), .A2(G141), .ZN(n702) );
  NAND2_X1 U776 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U777 ( .A1(G117), .A2(n878), .ZN(n704) );
  XNOR2_X1 U778 ( .A(KEYINPUT93), .B(n704), .ZN(n705) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n888) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n888), .ZN(n709) );
  XOR2_X1 U782 ( .A(KEYINPUT94), .B(n709), .Z(n718) );
  NAND2_X1 U783 ( .A1(G131), .A2(n882), .ZN(n711) );
  NAND2_X1 U784 ( .A1(G107), .A2(n878), .ZN(n710) );
  NAND2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U786 ( .A1(G95), .A2(n881), .ZN(n713) );
  NAND2_X1 U787 ( .A1(G119), .A2(n877), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U790 ( .A(n716), .B(KEYINPUT91), .ZN(n874) );
  AND2_X1 U791 ( .A1(n874), .A2(G1991), .ZN(n717) );
  NOR2_X1 U792 ( .A1(n718), .A2(n717), .ZN(n993) );
  INV_X1 U793 ( .A(n736), .ZN(n719) );
  NOR2_X1 U794 ( .A1(n993), .A2(n719), .ZN(n729) );
  INV_X1 U795 ( .A(n729), .ZN(n720) );
  NAND2_X1 U796 ( .A1(n733), .A2(n720), .ZN(n750) );
  INV_X1 U797 ( .A(n750), .ZN(n721) );
  AND2_X1 U798 ( .A1(n928), .A2(n721), .ZN(n722) );
  XNOR2_X1 U799 ( .A(G1986), .B(G290), .ZN(n917) );
  NAND2_X1 U800 ( .A1(n917), .A2(n736), .ZN(n738) );
  AND2_X1 U801 ( .A1(n722), .A2(n738), .ZN(n723) );
  NAND2_X1 U802 ( .A1(n724), .A2(n723), .ZN(n756) );
  AND2_X1 U803 ( .A1(n867), .A2(n725), .ZN(n726) );
  XNOR2_X1 U804 ( .A(n726), .B(KEYINPUT103), .ZN(n1008) );
  NOR2_X1 U805 ( .A1(G1996), .A2(n888), .ZN(n995) );
  NOR2_X1 U806 ( .A1(G1991), .A2(n874), .ZN(n990) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n727) );
  NOR2_X1 U808 ( .A1(n990), .A2(n727), .ZN(n728) );
  NOR2_X1 U809 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U810 ( .A1(n995), .A2(n730), .ZN(n731) );
  XNOR2_X1 U811 ( .A(KEYINPUT102), .B(n731), .ZN(n732) );
  XNOR2_X1 U812 ( .A(n732), .B(KEYINPUT39), .ZN(n734) );
  NAND2_X1 U813 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U814 ( .A1(n1008), .A2(n735), .ZN(n737) );
  NAND2_X1 U815 ( .A1(n737), .A2(n736), .ZN(n754) );
  INV_X1 U816 ( .A(n738), .ZN(n752) );
  NOR2_X1 U817 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XOR2_X1 U818 ( .A(n739), .B(KEYINPUT24), .Z(n740) );
  OR2_X1 U819 ( .A1(n745), .A2(n740), .ZN(n748) );
  NAND2_X1 U820 ( .A1(G8), .A2(G166), .ZN(n741) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n741), .ZN(n742) );
  XNOR2_X1 U822 ( .A(n742), .B(KEYINPUT101), .ZN(n744) );
  NAND2_X1 U823 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U824 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U825 ( .A1(n748), .A2(n747), .ZN(n749) );
  OR2_X1 U826 ( .A1(n750), .A2(n749), .ZN(n751) );
  OR2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U828 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U831 ( .A(G57), .ZN(G237) );
  INV_X1 U832 ( .A(G132), .ZN(G219) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  NAND2_X1 U834 ( .A1(G94), .A2(G452), .ZN(n758) );
  XNOR2_X1 U835 ( .A(n758), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U836 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U837 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U838 ( .A(G223), .ZN(n823) );
  NAND2_X1 U839 ( .A1(n823), .A2(G567), .ZN(n760) );
  XOR2_X1 U840 ( .A(KEYINPUT11), .B(n760), .Z(G234) );
  INV_X1 U841 ( .A(G860), .ZN(n766) );
  OR2_X1 U842 ( .A1(n934), .A2(n766), .ZN(G153) );
  INV_X1 U843 ( .A(G171), .ZN(G301) );
  INV_X1 U844 ( .A(G868), .ZN(n807) );
  NAND2_X1 U845 ( .A1(n920), .A2(n807), .ZN(n761) );
  XNOR2_X1 U846 ( .A(n761), .B(KEYINPUT74), .ZN(n763) );
  NAND2_X1 U847 ( .A1(G868), .A2(G301), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n763), .A2(n762), .ZN(G284) );
  NAND2_X1 U849 ( .A1(G868), .A2(G286), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G299), .A2(n807), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U852 ( .A1(n766), .A2(G559), .ZN(n767) );
  INV_X1 U853 ( .A(n920), .ZN(n794) );
  NAND2_X1 U854 ( .A1(n767), .A2(n794), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n934), .ZN(n769) );
  XOR2_X1 U857 ( .A(KEYINPUT79), .B(n769), .Z(n772) );
  NAND2_X1 U858 ( .A1(G868), .A2(n794), .ZN(n770) );
  NOR2_X1 U859 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U861 ( .A1(G123), .A2(n877), .ZN(n773) );
  XNOR2_X1 U862 ( .A(n773), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G99), .A2(n881), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT80), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G135), .A2(n882), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G111), .A2(n878), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n989) );
  XNOR2_X1 U870 ( .A(n989), .B(G2096), .ZN(n782) );
  INV_X1 U871 ( .A(G2100), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G67), .A2(n783), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G80), .A2(n784), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G93), .A2(n787), .ZN(n788) );
  XNOR2_X1 U877 ( .A(KEYINPUT81), .B(n788), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n791), .A2(G55), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n808) );
  NAND2_X1 U881 ( .A1(n794), .A2(G559), .ZN(n805) );
  XNOR2_X1 U882 ( .A(n934), .B(n805), .ZN(n795) );
  NOR2_X1 U883 ( .A1(G860), .A2(n795), .ZN(n796) );
  XOR2_X1 U884 ( .A(n808), .B(n796), .Z(G145) );
  XNOR2_X1 U885 ( .A(KEYINPUT19), .B(G305), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n797), .B(G288), .ZN(n798) );
  XNOR2_X1 U887 ( .A(KEYINPUT85), .B(n798), .ZN(n801) );
  XNOR2_X1 U888 ( .A(G290), .B(n799), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U890 ( .A(G166), .B(n802), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(n808), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n934), .B(n804), .ZN(n895) );
  XNOR2_X1 U893 ( .A(n805), .B(n895), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n806), .A2(G868), .ZN(n810) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U897 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U903 ( .A1(G220), .A2(G219), .ZN(n815) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(n815), .Z(n816) );
  NOR2_X1 U905 ( .A1(G218), .A2(n816), .ZN(n817) );
  NAND2_X1 U906 ( .A1(G96), .A2(n817), .ZN(n827) );
  NAND2_X1 U907 ( .A1(n827), .A2(G2106), .ZN(n821) );
  NAND2_X1 U908 ( .A1(G120), .A2(G108), .ZN(n818) );
  NOR2_X1 U909 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U910 ( .A1(G69), .A2(n819), .ZN(n828) );
  NAND2_X1 U911 ( .A1(n828), .A2(G567), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n830) );
  NAND2_X1 U913 ( .A1(G661), .A2(G483), .ZN(n822) );
  NOR2_X1 U914 ( .A1(n830), .A2(n822), .ZN(n826) );
  NAND2_X1 U915 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT105), .B(n829), .Z(G325) );
  XOR2_X1 U925 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(n830), .ZN(G319) );
  XOR2_X1 U929 ( .A(G2100), .B(KEYINPUT108), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2678), .B(KEYINPUT43), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2090), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U936 ( .A(KEYINPUT107), .B(G2096), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U938 ( .A(G2078), .B(G2084), .Z(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U943 ( .A(G1981), .B(G1956), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(n849), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G124), .A2(n877), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n852), .B(KEYINPUT44), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT110), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G100), .A2(n881), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G136), .A2(n882), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G112), .A2(n878), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G103), .A2(n881), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G139), .A2(n882), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n877), .A2(G127), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G115), .A2(n878), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(KEYINPUT47), .B(n864), .Z(n865) );
  NOR2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n1001) );
  XOR2_X1 U968 ( .A(G162), .B(n1001), .Z(n869) );
  XOR2_X1 U969 ( .A(G164), .B(n867), .Z(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n873), .B(n872), .Z(n876) );
  XOR2_X1 U975 ( .A(n874), .B(n989), .Z(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n892) );
  NAND2_X1 U977 ( .A1(n877), .A2(G130), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U980 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U986 ( .A(G160), .B(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U988 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U989 ( .A(G171), .B(n920), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(G286), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2438), .B(KEYINPUT104), .Z(n899) );
  XNOR2_X1 U994 ( .A(G2443), .B(G2430), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(n900), .B(G2435), .Z(n902) );
  XNOR2_X1 U997 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U999 ( .A(G2451), .B(G2427), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G2454), .B(G2446), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1002 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1003 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  INV_X1 U1012 ( .A(n913), .ZN(G401) );
  NAND2_X1 U1013 ( .A1(G1971), .A2(G303), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n926) );
  XNOR2_X1 U1015 ( .A(G1956), .B(G299), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n924) );
  XNOR2_X1 U1017 ( .A(G171), .B(G1961), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(G1348), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT121), .B(n927), .Z(n933) );
  XNOR2_X1 U1024 ( .A(G168), .B(G1966), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n930), .B(KEYINPUT57), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT120), .B(n931), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G1341), .B(n934), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1031 ( .A(KEYINPUT122), .B(n937), .Z(n939) );
  XNOR2_X1 U1032 ( .A(G16), .B(KEYINPUT56), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n1021) );
  XNOR2_X1 U1034 ( .A(G5), .B(G1961), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(KEYINPUT123), .ZN(n960) );
  XNOR2_X1 U1036 ( .A(n941), .B(G20), .ZN(n949) );
  XOR2_X1 U1037 ( .A(G1981), .B(G6), .Z(n944) );
  XOR2_X1 U1038 ( .A(G19), .B(KEYINPUT124), .Z(n942) );
  XNOR2_X1 U1039 ( .A(G1341), .B(n942), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1041 ( .A(KEYINPUT59), .B(G1348), .Z(n945) );
  XNOR2_X1 U1042 ( .A(G4), .B(n945), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(n950), .B(KEYINPUT60), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G22), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G23), .B(G1976), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G1986), .B(KEYINPUT125), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n953), .B(G24), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(G21), .B(G1966), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n963), .Z(n964) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n964), .ZN(n965) );
  XOR2_X1 U1059 ( .A(KEYINPUT126), .B(n965), .Z(n966) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n966), .ZN(n1019) );
  XOR2_X1 U1061 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT54), .B(n967), .ZN(n984) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n982) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n978) );
  XOR2_X1 U1067 ( .A(G25), .B(G1991), .Z(n970) );
  NAND2_X1 U1068 ( .A1(n970), .A2(G28), .ZN(n976) );
  XOR2_X1 U1069 ( .A(G1996), .B(G32), .Z(n973) );
  XNOR2_X1 U1070 ( .A(n971), .B(G27), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(KEYINPUT116), .B(n974), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n980), .B(KEYINPUT117), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n985), .B(KEYINPUT118), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT55), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(G29), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n988), .B(KEYINPUT119), .ZN(n1017) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(KEYINPUT114), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n1011) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n996), .Z(n1000) );
  XOR2_X1 U1089 ( .A(G160), .B(G2084), .Z(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G2072), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G164), .B(G2078), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT115), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(KEYINPUT52), .ZN(n1014) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(G29), .A2(n1015), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

