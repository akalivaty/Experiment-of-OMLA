//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT71), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(KEYINPUT71), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  AND2_X1   g041(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G101), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT74), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n477), .A2(new_n474), .A3(G101), .A4(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT3), .B1(new_n480), .B2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(G137), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n479), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n490));
  INV_X1    g065(.A(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT73), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(G137), .A3(new_n469), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT75), .A3(new_n479), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n473), .B1(new_n489), .B2(new_n496), .ZN(G160));
  NOR2_X1   g072(.A1(new_n483), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G136), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n483), .A2(new_n469), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G124), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT77), .ZN(new_n504));
  OAI221_X1 g079(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n506), .B(new_n507), .ZN(G162));
  NAND3_X1  g083(.A1(new_n484), .A2(G138), .A3(new_n485), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT4), .B1(new_n483), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n490), .A2(G2104), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G138), .ZN(new_n515));
  NOR3_X1   g090(.A1(new_n467), .A2(new_n468), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(KEYINPUT79), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT79), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n510), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n494), .A2(G126), .A3(G2105), .ZN(new_n522));
  OR2_X1    g097(.A1(G102), .A2(G2105), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n523), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n521), .A2(KEYINPUT80), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT80), .B1(new_n521), .B2(new_n526), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(G164));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G50), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT5), .B(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n538), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n532), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G166));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n547));
  AOI22_X1  g122(.A1(G51), .A2(new_n535), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT5), .B(G543), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n537), .A2(G89), .ZN(new_n551));
  NAND2_X1  g126(.A1(G63), .A2(G651), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n549), .A2(new_n553), .ZN(G168));
  AOI22_X1  g129(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n532), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n535), .A2(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n539), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n559), .A2(KEYINPUT81), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(KEYINPUT81), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  NAND2_X1  g138(.A1(new_n535), .A2(G43), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT82), .B(G81), .Z(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n539), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n532), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g146(.A(KEYINPUT83), .B(KEYINPUT8), .Z(new_n572));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n539), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT84), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n535), .A2(G53), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT9), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n538), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n532), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(G299));
  INV_X1    g160(.A(G168), .ZN(G286));
  INV_X1    g161(.A(G166), .ZN(G303));
  NAND2_X1  g162(.A1(new_n579), .A2(G87), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n538), .A2(G74), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G49), .B2(new_n535), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n550), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G48), .B2(new_n535), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n577), .A2(new_n578), .A3(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT85), .ZN(G305));
  INV_X1    g173(.A(new_n539), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G85), .B1(G47), .B2(new_n535), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT87), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n532), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT86), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n535), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n538), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n532), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n579), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n577), .A2(new_n578), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n609), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  XNOR2_X1  g195(.A(G280), .B(KEYINPUT88), .ZN(G297));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g201(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n627));
  XNOR2_X1  g202(.A(G323), .B(new_n627), .ZN(G282));
  NOR2_X1   g203(.A1(new_n491), .A2(G2105), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n470), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(G2100), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n632), .B2(new_n631), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n635), .A2(new_n633), .A3(G2100), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n633), .B2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n498), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n502), .A2(G123), .ZN(new_n639));
  OAI221_X1 g214(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT91), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT92), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT93), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n666), .B1(new_n663), .B2(new_n665), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n678), .A2(new_n683), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n686));
  AOI211_X1 g261(.A(new_n682), .B(new_n684), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1981), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT98), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT99), .Z(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G1971), .ZN(new_n706));
  MUX2_X1   g281(.A(G23), .B(G288), .S(G16), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(G1971), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n701), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  MUX2_X1   g290(.A(G24), .B(G290), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(new_n695), .ZN(new_n717));
  AOI22_X1  g292(.A1(G119), .A2(new_n502), .B1(new_n498), .B2(G131), .ZN(new_n718));
  NOR2_X1   g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT97), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G25), .B(new_n722), .S(G29), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT36), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n728), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT29), .Z(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT103), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n728), .A2(G32), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n498), .A2(G141), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n502), .A2(G129), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT26), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n740), .A2(new_n741), .B1(G105), .B2(new_n629), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n736), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n735), .B1(new_n744), .B2(new_n728), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n728), .A2(G33), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  INV_X1    g325(.A(new_n469), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n470), .A2(G127), .ZN(new_n752));
  INV_X1    g327(.A(G115), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n491), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n751), .A2(new_n754), .B1(new_n498), .B2(G139), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n748), .B1(new_n756), .B2(new_n728), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n747), .B1(G2072), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n760), .B2(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(KEYINPUT24), .B2(new_n760), .ZN(new_n762));
  INV_X1    g337(.A(G160), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n728), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n758), .B1(G2072), .B2(new_n757), .C1(new_n759), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT101), .ZN(new_n766));
  NOR2_X1   g341(.A1(G286), .A2(new_n702), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT102), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT102), .B1(G16), .B2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n771), .A2(G1966), .B1(new_n745), .B2(new_n746), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G1966), .B2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n728), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT28), .Z(new_n775));
  OAI221_X1 g350(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(G128), .A2(new_n502), .B1(new_n498), .B2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n764), .A2(new_n759), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n702), .A2(G5), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G171), .B2(new_n702), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G1961), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G28), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT30), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(KEYINPUT30), .ZN(new_n790));
  OR2_X1    g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n789), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n641), .B2(new_n728), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n569), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G16), .B2(G19), .ZN(new_n796));
  INV_X1    g371(.A(G1341), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n798), .B1(new_n797), .B2(new_n796), .C1(new_n785), .C2(G1961), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n773), .A2(new_n787), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n702), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n619), .B2(new_n702), .ZN(new_n803));
  INV_X1    g378(.A(G1956), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n615), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1348), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n728), .A2(G27), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G164), .B2(new_n728), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n800), .A2(new_n805), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  AOI211_X1 g389(.A(new_n766), .B(new_n814), .C1(new_n731), .C2(new_n732), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n727), .A2(new_n734), .A3(new_n815), .ZN(G311));
  NAND3_X1  g391(.A1(new_n727), .A2(new_n734), .A3(new_n815), .ZN(G150));
  NAND2_X1  g392(.A1(new_n535), .A2(G55), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n539), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n532), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n615), .A2(G559), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT38), .Z(new_n828));
  INV_X1    g403(.A(new_n823), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT104), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n569), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n569), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n828), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n824), .B1(new_n839), .B2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n826), .B1(new_n840), .B2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(KEYINPUT107), .B(G37), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(new_n763), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n641), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT105), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n756), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n744), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n498), .A2(G142), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n502), .A2(G130), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n631), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n849), .B(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT79), .B1(new_n514), .B2(new_n516), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n513), .B1(new_n516), .B2(new_n494), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n525), .B1(new_n858), .B2(new_n517), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n780), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n722), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n855), .B(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n844), .B1(new_n846), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n846), .ZN(new_n864));
  INV_X1    g439(.A(new_n862), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT106), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT106), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g444(.A1(new_n829), .A2(G868), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n624), .B(KEYINPUT108), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n837), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n615), .A2(KEYINPUT109), .A3(G299), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT109), .B1(new_n615), .B2(G299), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n615), .A2(G299), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n873), .A2(new_n874), .A3(new_n878), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n872), .A2(new_n876), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT110), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(G305), .A2(G290), .ZN(new_n884));
  NAND2_X1  g459(.A1(G305), .A2(G290), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G288), .B(G303), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n887), .A3(new_n885), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT110), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n870), .B1(new_n895), .B2(G868), .ZN(G295));
  AOI21_X1  g471(.A(new_n870), .B1(new_n895), .B2(G868), .ZN(G331));
  NAND2_X1  g472(.A1(G301), .A2(G168), .ZN(new_n898));
  OAI211_X1 g473(.A(G286), .B(new_n556), .C1(new_n561), .C2(new_n560), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n836), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n569), .B1(new_n830), .B2(new_n832), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n835), .A2(new_n836), .A3(new_n899), .A4(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n877), .A2(new_n905), .A3(new_n879), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n876), .A2(new_n903), .A3(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n891), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n891), .A3(new_n907), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n844), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT111), .B1(new_n912), .B2(new_n913), .ZN(new_n919));
  INV_X1    g494(.A(new_n911), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n891), .B1(new_n906), .B2(new_n907), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n843), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n917), .B1(new_n915), .B2(new_n913), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n925), .A2(KEYINPUT112), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT112), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(G397));
  INV_X1    g504(.A(G2067), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n780), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT113), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n744), .ZN(new_n933));
  INV_X1    g508(.A(new_n473), .ZN(new_n934));
  INV_X1    g509(.A(new_n496), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT75), .B1(new_n495), .B2(new_n479), .ZN(new_n936));
  OAI211_X1 g511(.A(G40), .B(new_n934), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G1384), .B1(new_n521), .B2(new_n526), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT45), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n941), .A3(new_n744), .ZN(new_n944));
  INV_X1    g519(.A(new_n724), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n722), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G2067), .B2(new_n780), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n939), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n943), .A2(new_n944), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n722), .A2(new_n945), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n939), .B1(new_n951), .B2(new_n946), .ZN(new_n952));
  NOR2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n939), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT48), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n933), .A2(new_n939), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT126), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n939), .A2(new_n941), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(KEYINPUT125), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(new_n960), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT47), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n957), .A2(new_n968), .A3(new_n960), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n949), .A2(new_n956), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n972), .B(new_n973), .C1(new_n527), .C2(new_n528), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n521), .A2(new_n526), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n973), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n937), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n804), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n619), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(G299), .A2(KEYINPUT117), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(G1384), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n937), .B1(new_n975), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT56), .B(G2072), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT80), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n975), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n521), .A2(KEYINPUT80), .A3(new_n526), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n988), .B(new_n989), .C1(new_n993), .C2(KEYINPUT45), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n979), .A2(new_n985), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n938), .A2(new_n972), .ZN(new_n996));
  INV_X1    g571(.A(new_n937), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n996), .B(new_n997), .C1(new_n993), .C2(new_n972), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n976), .A2(new_n937), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n998), .A2(new_n808), .B1(new_n930), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n615), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n985), .B1(new_n979), .B2(new_n994), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT61), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n979), .A2(new_n985), .A3(new_n994), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(new_n1003), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(G1341), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n976), .B2(new_n937), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n987), .ZN(new_n1012));
  OAI211_X1 g587(.A(G40), .B(G160), .C1(new_n859), .C2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n973), .B1(new_n527), .B2(new_n528), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(new_n986), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1015), .B2(new_n941), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n569), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT59), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n941), .B(new_n988), .C1(new_n993), .C2(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n1010), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n1017), .A3(new_n1022), .A4(new_n569), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n983), .A2(new_n984), .ZN(new_n1025));
  INV_X1    g600(.A(new_n994), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1956), .B1(new_n974), .B2(new_n977), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT61), .A3(new_n995), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1000), .A2(KEYINPUT60), .A3(new_n1001), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1007), .A2(new_n1024), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1000), .A2(KEYINPUT60), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1000), .A2(KEYINPUT60), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n1001), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1004), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n859), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(new_n732), .A3(new_n997), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n988), .B1(new_n993), .B2(KEYINPUT45), .ZN(new_n1040));
  INV_X1    g615(.A(G1971), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1036), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G166), .A2(new_n1036), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  OAI22_X1  g622(.A1(G166), .A2(new_n1036), .B1(KEYINPUT114), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1015), .A2(G1971), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n978), .A2(G2090), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1049), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT115), .B1(new_n597), .B2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n595), .A2(new_n596), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n599), .A2(G86), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n595), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1063), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n999), .A2(new_n1036), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n588), .A2(G1976), .A3(new_n590), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1069), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1050), .A2(new_n1055), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1040), .B2(G2078), .ZN(new_n1079));
  INV_X1    g654(.A(G1961), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n998), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n937), .B1(new_n976), .B2(new_n986), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n987), .B1(new_n527), .B2(new_n528), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT53), .A4(new_n812), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  OAI211_X1 g662(.A(G40), .B(G160), .C1(new_n938), .C2(KEYINPUT45), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT53), .B(new_n812), .C1(new_n859), .C2(new_n1012), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1079), .B(new_n1081), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1090), .B2(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1077), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n937), .A2(G2084), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1094));
  INV_X1    g669(.A(G1966), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1038), .A2(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G168), .A2(new_n1036), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT51), .B1(new_n1097), .B2(KEYINPUT121), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1098), .B(new_n1100), .C1(new_n1096), .C2(new_n1036), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1100), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n996), .B(new_n1093), .C1(new_n993), .C2(new_n972), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1012), .B1(new_n991), .B2(new_n992), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1095), .B1(new_n1104), .B2(new_n1088), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(G8), .B(new_n1102), .C1(new_n1106), .C2(G286), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1099), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1085), .A2(G171), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(G171), .B2(new_n1090), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1035), .A2(new_n1092), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT123), .B(KEYINPUT62), .C1(new_n1114), .C2(new_n1099), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1077), .A2(new_n1109), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1076), .A2(new_n1049), .A3(new_n1043), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1060), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G288), .A2(G1976), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1069), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1068), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g702(.A(KEYINPUT116), .B(new_n1123), .C1(new_n1069), .C2(new_n1124), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1106), .A2(G8), .A3(G168), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1077), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1130), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1133), .A2(new_n1050), .A3(new_n1076), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1129), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1113), .A2(new_n1121), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n695), .B1(new_n601), .B2(new_n604), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n939), .B1(new_n953), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n950), .A2(new_n1139), .A3(new_n952), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1137), .A2(KEYINPUT124), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT124), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n971), .B1(new_n1141), .B2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g718(.A1(G401), .A2(G229), .A3(new_n465), .A4(G227), .ZN(new_n1145));
  NAND3_X1  g719(.A1(new_n1145), .A2(new_n868), .A3(new_n916), .ZN(G225));
  INV_X1    g720(.A(G225), .ZN(G308));
endmodule


