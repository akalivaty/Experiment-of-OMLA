//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT68), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(KEYINPUT23), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT25), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n206), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n220), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n207), .A4(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n225), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n211), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n213), .A2(new_n214), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT64), .Z(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT33), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n205), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(KEYINPUT32), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n240), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n241), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n250));
  NOR2_X1   g049(.A1(new_n242), .A2(KEYINPUT34), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n249), .A2(new_n250), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n243), .B(KEYINPUT32), .C1(new_n244), .C2(new_n205), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n247), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT36), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT83), .B(G155gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(G162gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT84), .ZN(new_n261));
  XOR2_X1   g060(.A(G155gat), .B(G162gat), .Z(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G148gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT82), .ZN(new_n265));
  INV_X1    g064(.A(G148gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G141gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(KEYINPUT82), .A3(G141gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G155gat), .ZN(new_n271));
  INV_X1    g070(.A(G162gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT2), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n273), .A2(new_n274), .B1(new_n264), .B2(new_n267), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n274), .B2(new_n273), .ZN(new_n276));
  XNOR2_X1  g075(.A(G155gat), .B(G162gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n261), .A2(new_n270), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n285), .B(new_n258), .C1(new_n259), .C2(G162gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n270), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(new_n279), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT85), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT29), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  XNOR2_X1  g094(.A(G197gat), .B(G204gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT70), .B(G218gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT22), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT72), .B1(new_n301), .B2(KEYINPUT71), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n292), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n291), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT86), .B1(new_n301), .B2(new_n292), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n301), .A2(new_n292), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n301), .A2(KEYINPUT86), .A3(new_n292), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n289), .B1(new_n311), .B2(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT31), .B(G50gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G22gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n299), .A2(new_n300), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT71), .A3(new_n296), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n292), .B1(new_n323), .B2(new_n293), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n295), .A2(new_n301), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n302), .B(KEYINPUT73), .C1(new_n292), .C2(new_n303), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n291), .A2(KEYINPUT88), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT88), .ZN(new_n331));
  AOI211_X1 g130(.A(new_n331), .B(KEYINPUT29), .C1(new_n283), .C2(new_n290), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n282), .B1(new_n304), .B2(KEYINPUT29), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n334), .A2(KEYINPUT87), .A3(new_n289), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT87), .B1(new_n334), .B2(new_n289), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n316), .B(new_n320), .C1(new_n339), .C2(new_n313), .ZN(new_n340));
  INV_X1    g139(.A(new_n320), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n313), .B1(new_n333), .B2(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(new_n315), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n238), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n289), .A2(KEYINPUT85), .A3(KEYINPUT3), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n287), .A2(new_n288), .A3(new_n238), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT4), .A4(new_n238), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n289), .B(new_n238), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(new_n349), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT5), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT0), .ZN(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT90), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n356), .B2(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n283), .A2(new_n290), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n354), .B1(new_n372), .B2(new_n345), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT5), .B1(new_n373), .B2(new_n349), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n365), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n358), .B1(new_n373), .B2(new_n349), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n366), .B(new_n368), .C1(new_n376), .C2(new_n367), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n371), .A2(new_n374), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT90), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT6), .A4(new_n366), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n370), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT77), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT78), .Z(new_n388));
  INV_X1    g187(.A(KEYINPUT38), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n234), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n217), .A2(KEYINPUT25), .B1(new_n231), .B2(new_n232), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n394), .B2(new_n230), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n395), .B2(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n304), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n329), .B2(new_n396), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n390), .B1(new_n398), .B2(KEYINPUT37), .ZN(new_n399));
  INV_X1    g198(.A(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n305), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n329), .A2(new_n396), .A3(KEYINPUT75), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT75), .B1(new_n329), .B2(new_n396), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n404), .B2(KEYINPUT37), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n400), .B2(new_n328), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n329), .A2(new_n396), .A3(KEYINPUT75), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n407), .A2(new_n408), .B1(new_n305), .B2(new_n400), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n387), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n401), .C1(new_n402), .C2(new_n403), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(KEYINPUT37), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n387), .B1(new_n409), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(new_n418), .B2(KEYINPUT38), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n383), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n412), .A2(new_n414), .A3(new_n388), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n409), .A2(KEYINPUT30), .A3(new_n387), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT40), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT89), .B1(new_n373), .B2(new_n349), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n348), .A2(new_n355), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n429));
  INV_X1    g228(.A(new_n349), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n357), .B2(new_n349), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n365), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT39), .B1(new_n427), .B2(new_n431), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n426), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(KEYINPUT40), .A3(new_n365), .A4(new_n434), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n425), .A2(new_n437), .A3(new_n439), .A4(new_n377), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n344), .B1(new_n420), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n424), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n442), .A2(new_n443), .B1(new_n422), .B2(new_n410), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n421), .A2(KEYINPUT79), .A3(new_n424), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n379), .A2(new_n369), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n344), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n257), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n340), .A2(new_n343), .A3(new_n256), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n340), .A2(new_n343), .A3(new_n256), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n453), .A2(KEYINPUT35), .A3(new_n425), .ZN(new_n454));
  INV_X1    g253(.A(new_n383), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n449), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G183gat), .B(G211gat), .Z(new_n458));
  INV_X1    g257(.A(KEYINPUT95), .ZN(new_n459));
  INV_X1    g258(.A(G57gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(G64gat), .ZN(new_n461));
  INV_X1    g260(.A(G64gat), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT95), .B1(new_n462), .B2(G57gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(G57gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G71gat), .A2(G78gat), .ZN(new_n466));
  OR2_X1    g265(.A1(G71gat), .A2(G78gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n466), .B(new_n467), .C1(new_n471), .C2(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT21), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G231gat), .A2(G233gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G127gat), .B(G155gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT96), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n479), .B(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  INV_X1    g282(.A(G1gat), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n484), .A2(KEYINPUT16), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(new_n484), .ZN(new_n487));
  OAI21_X1  g286(.A(G8gat), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n485), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n489), .B(new_n490), .C1(new_n484), .C2(new_n483), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n474), .B2(new_n473), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n482), .A2(new_n493), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n458), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n482), .A2(new_n493), .ZN(new_n498));
  INV_X1    g297(.A(new_n458), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(G232gat), .A2(G233gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(KEYINPUT41), .ZN(new_n503));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  OR3_X1    g304(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n506), .A2(new_n507), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT91), .B1(new_n510), .B2(G50gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  INV_X1    g311(.A(G50gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(G43gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT92), .B(G50gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(G43gat), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n510), .B2(G50gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n510), .B2(G50gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n509), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n509), .A2(new_n521), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT8), .ZN(new_n527));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G85gat), .ZN(new_n531));
  INV_X1    g330(.A(G92gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n527), .A2(new_n530), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G99gat), .B(G106gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(KEYINPUT98), .A3(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(KEYINPUT8), .A2(new_n526), .B1(new_n531), .B2(new_n532), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n539), .A2(new_n536), .A3(new_n530), .A4(new_n534), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT98), .B1(new_n535), .B2(new_n537), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n525), .A2(new_n543), .B1(KEYINPUT41), .B2(new_n502), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT92), .B(G50gat), .Z(new_n545));
  AOI22_X1  g344(.A1(new_n545), .A2(new_n510), .B1(new_n511), .B2(new_n514), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n521), .B1(new_n546), .B2(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n508), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n523), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT17), .B1(new_n522), .B2(new_n524), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n552), .B2(new_n543), .ZN(new_n553));
  XOR2_X1   g352(.A(G190gat), .B(G218gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n505), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n557), .B(new_n559), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n501), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n488), .A2(new_n491), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n488), .B2(new_n491), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n551), .A3(new_n550), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n565), .A2(new_n550), .A3(new_n551), .A4(KEYINPUT94), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n525), .A2(new_n488), .A3(new_n491), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n570), .A2(new_n571), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n569), .A4(new_n568), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n525), .B(new_n492), .Z(new_n577));
  XOR2_X1   g376(.A(new_n569), .B(KEYINPUT13), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT11), .ZN(new_n582));
  INV_X1    g381(.A(G169gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT12), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n574), .A2(new_n576), .A3(new_n579), .A4(new_n586), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n473), .B1(new_n541), .B2(new_n542), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n535), .A2(new_n537), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(new_n470), .A3(new_n472), .A4(new_n540), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT100), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n460), .A2(G64gat), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT9), .B1(new_n464), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n467), .A2(new_n466), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n465), .A2(new_n469), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n593), .A4(new_n540), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n592), .A2(new_n595), .A3(new_n596), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n543), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n603), .A2(KEYINPUT101), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT101), .B1(new_n603), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n591), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT102), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n609), .B(new_n591), .C1(new_n605), .C2(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n595), .A3(new_n602), .ZN(new_n612));
  INV_X1    g411(.A(new_n591), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT103), .B1(new_n620), .B2(new_n591), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n622), .B(new_n613), .C1(new_n603), .C2(new_n604), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n617), .B1(new_n624), .B2(new_n614), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n561), .A2(new_n590), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n457), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n446), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n425), .ZN(new_n632));
  NOR2_X1   g431(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n632), .A2(G8gat), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(G8gat), .B1(new_n632), .B2(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(new_n632), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n635), .B(new_n636), .C1(KEYINPUT42), .C2(new_n637), .ZN(G1325gat));
  AOI21_X1  g437(.A(G15gat), .B1(new_n628), .B2(new_n256), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT105), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(KEYINPUT105), .ZN(new_n641));
  INV_X1    g440(.A(new_n257), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G15gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT106), .Z(new_n644));
  AOI22_X1  g443(.A1(new_n640), .A2(new_n641), .B1(new_n628), .B2(new_n644), .ZN(G1326gat));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n344), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT107), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT43), .B(G22gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  XNOR2_X1  g448(.A(new_n557), .B(new_n559), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n501), .A2(new_n590), .A3(new_n626), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n457), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n446), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT45), .Z(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n451), .A2(KEYINPUT35), .B1(new_n454), .B2(new_n455), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n425), .A2(new_n377), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n437), .A2(new_n439), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n657), .A2(new_n658), .B1(new_n383), .B2(new_n419), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n447), .B1(new_n659), .B2(new_n344), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n660), .B2(new_n257), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n655), .B1(new_n661), .B2(new_n560), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n420), .A2(new_n440), .ZN(new_n663));
  INV_X1    g462(.A(new_n344), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n642), .B1(new_n665), .B2(new_n447), .ZN(new_n666));
  OAI211_X1 g465(.A(KEYINPUT44), .B(new_n650), .C1(new_n666), .C2(new_n656), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n651), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668), .B2(new_n446), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n669), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671));
  INV_X1    g470(.A(G36gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n425), .A2(new_n672), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n652), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n652), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n425), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n668), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT108), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n676), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1329gat));
  INV_X1    g482(.A(new_n256), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n510), .B1(new_n652), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n642), .A2(G43gat), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n668), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g487(.A(new_n545), .B1(new_n668), .B2(new_n664), .ZN(new_n689));
  INV_X1    g488(.A(new_n652), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n344), .A3(new_n516), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT48), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n692), .B(new_n694), .ZN(G1331gat));
  NAND2_X1  g494(.A1(new_n588), .A2(new_n589), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n561), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n457), .A2(new_n626), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n629), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT110), .B(G57gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1332gat));
  INV_X1    g500(.A(KEYINPUT49), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n698), .B(new_n425), .C1(new_n702), .C2(new_n462), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n462), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1333gat));
  NAND2_X1  g504(.A1(new_n698), .A2(new_n642), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n684), .A2(G71gat), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n706), .A2(G71gat), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g508(.A1(new_n698), .A2(new_n344), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  INV_X1    g510(.A(new_n501), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n590), .ZN(new_n713));
  INV_X1    g512(.A(new_n626), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT111), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n662), .A2(new_n667), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n662), .A2(new_n667), .A3(KEYINPUT112), .A4(new_n716), .ZN(new_n720));
  AND4_X1   g519(.A1(G85gat), .A2(new_n719), .A3(new_n629), .A4(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n713), .B1(KEYINPUT113), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n457), .A2(new_n650), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(KEYINPUT113), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n457), .A2(new_n650), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n726), .A2(new_n629), .A3(new_n626), .A4(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n721), .B1(new_n531), .B2(new_n729), .ZN(G1336gat));
  OAI21_X1  g529(.A(G92gat), .B1(new_n717), .B2(new_n677), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n677), .A2(G92gat), .A3(new_n714), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n726), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n733), .B(KEYINPUT114), .Z(new_n736));
  AND3_X1   g535(.A1(new_n726), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n425), .A3(new_n720), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(G92gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(new_n732), .ZN(G1337gat));
  AND4_X1   g539(.A1(G99gat), .A2(new_n719), .A3(new_n642), .A4(new_n720), .ZN(new_n741));
  INV_X1    g540(.A(G99gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n256), .A3(new_n626), .A4(new_n728), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(G1338gat));
  OAI21_X1  g543(.A(G106gat), .B1(new_n717), .B2(new_n664), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n664), .A2(G106gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n626), .A3(new_n728), .A4(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AND4_X1   g548(.A1(new_n626), .A2(new_n726), .A3(new_n728), .A4(new_n746), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n719), .A2(new_n344), .A3(new_n720), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G106gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n752), .B2(new_n748), .ZN(G1339gat));
  NOR3_X1   g552(.A1(new_n561), .A2(new_n696), .A3(new_n626), .ZN(new_n754));
  INV_X1    g553(.A(new_n619), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n603), .A2(new_n613), .A3(new_n604), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT54), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n620), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n603), .A2(KEYINPUT101), .A3(new_n604), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n609), .B1(new_n762), .B2(new_n591), .ZN(new_n763));
  INV_X1    g562(.A(new_n610), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n621), .B2(new_n623), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n617), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(KEYINPUT55), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n617), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n611), .B2(new_n758), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n755), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n569), .B1(new_n575), .B2(new_n568), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n577), .A2(new_n578), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n585), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n589), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n765), .A2(new_n768), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n775), .A2(new_n650), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n626), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n782), .A2(new_n696), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n787), .B2(new_n650), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n754), .B1(new_n788), .B2(new_n712), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n446), .A2(new_n425), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n453), .ZN(new_n793));
  AOI21_X1  g592(.A(G113gat), .B1(new_n793), .B2(new_n696), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n793), .B(KEYINPUT116), .Z(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n696), .A2(G113gat), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G1340gat));
  AOI21_X1  g597(.A(G120gat), .B1(new_n793), .B2(new_n626), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n626), .A2(G120gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n796), .B2(new_n800), .ZN(G1341gat));
  OAI21_X1  g600(.A(G127gat), .B1(new_n795), .B2(new_n712), .ZN(new_n802));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n793), .A2(new_n803), .A3(new_n501), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1342gat));
  OAI21_X1  g604(.A(G134gat), .B1(new_n795), .B2(new_n560), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n560), .A2(new_n425), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT117), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(G134gat), .A3(new_n453), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n790), .A3(new_n629), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT56), .Z(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n811), .ZN(G1343gat));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT115), .B1(new_n773), .B2(KEYINPUT55), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n757), .B1(new_n608), .B2(new_n610), .ZN(new_n815));
  NOR4_X1   g614(.A1(new_n815), .A2(new_n772), .A3(new_n770), .A4(new_n781), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n619), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n782), .A2(new_n696), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n784), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n560), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n501), .B1(new_n820), .B2(new_n783), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n813), .B(new_n344), .C1(new_n821), .C2(new_n754), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n791), .A2(new_n257), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n765), .A2(new_n827), .A3(new_n768), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT118), .B1(new_n815), .B2(new_n772), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n781), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n696), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n784), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n832), .A2(KEYINPUT119), .A3(new_n560), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT119), .B1(new_n832), .B2(new_n560), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n783), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n712), .ZN(new_n836));
  INV_X1    g635(.A(new_n754), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n664), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n826), .B1(new_n838), .B2(new_n813), .ZN(new_n839));
  OAI21_X1  g638(.A(G141gat), .B1(new_n839), .B2(new_n590), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n642), .A2(new_n664), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n792), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n696), .A2(new_n263), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT120), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n783), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(new_n780), .B2(KEYINPUT118), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n590), .B1(new_n852), .B2(new_n828), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n785), .B1(new_n853), .B2(new_n775), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n854), .B2(new_n650), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n832), .A2(KEYINPUT119), .A3(new_n560), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n837), .B1(new_n857), .B2(new_n501), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n344), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n825), .B1(new_n859), .B2(KEYINPUT57), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n263), .B1(new_n860), .B2(new_n696), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n848), .A2(new_n841), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT58), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n849), .A2(new_n863), .ZN(G1344gat));
  XOR2_X1   g663(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n865));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n789), .B2(new_n664), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n664), .A2(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n832), .A2(new_n560), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n501), .B1(new_n868), .B2(new_n783), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n869), .B2(new_n754), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n866), .A2(new_n626), .A3(new_n870), .A4(new_n824), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n865), .B1(new_n871), .B2(G148gat), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n826), .B(new_n626), .C1(new_n838), .C2(new_n813), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n266), .A2(KEYINPUT59), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n789), .A2(new_n446), .A3(new_n844), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n876), .A2(new_n266), .A3(new_n677), .A4(new_n626), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT123), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(new_n874), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n860), .B2(new_n626), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n877), .C1(new_n882), .C2(new_n872), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n883), .ZN(G1345gat));
  AOI21_X1  g683(.A(new_n259), .B1(new_n845), .B2(new_n501), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n501), .A2(new_n259), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n860), .B2(new_n886), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n839), .B2(new_n560), .ZN(new_n888));
  INV_X1    g687(.A(new_n808), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n876), .A2(new_n272), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1347gat));
  NAND2_X1  g690(.A1(new_n446), .A2(new_n425), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n789), .A2(new_n453), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n696), .ZN(new_n894));
  INV_X1    g693(.A(new_n892), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT124), .B1(new_n895), .B2(new_n256), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n892), .A2(new_n897), .A3(new_n684), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n896), .A2(new_n344), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n790), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT125), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n790), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n590), .A2(new_n583), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(G1348gat));
  OAI21_X1  g706(.A(G176gat), .B1(new_n904), .B2(new_n714), .ZN(new_n908));
  INV_X1    g707(.A(G176gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n909), .A3(new_n626), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1349gat));
  AND2_X1   g710(.A1(new_n501), .A2(new_n225), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT126), .B1(new_n893), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n904), .A2(new_n712), .ZN(new_n914));
  INV_X1    g713(.A(G183gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n918), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n893), .A2(new_n227), .A3(new_n650), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n650), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(G190gat), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT61), .B(new_n227), .C1(new_n905), .C2(new_n650), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  NOR3_X1   g725(.A1(new_n789), .A2(new_n844), .A3(new_n892), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n696), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n257), .A2(new_n866), .A3(new_n870), .A4(new_n895), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n696), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(new_n927), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(G204gat), .A3(new_n714), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n866), .A2(new_n626), .A3(new_n870), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n895), .A2(new_n257), .ZN(new_n936));
  OAI21_X1  g735(.A(G204gat), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1353gat));
  OR3_X1    g737(.A1(new_n932), .A2(G211gat), .A3(new_n712), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n929), .A2(new_n501), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n927), .B2(new_n650), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT127), .Z(new_n945));
  AND2_X1   g744(.A1(new_n650), .A2(new_n298), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1355gat));
endmodule


