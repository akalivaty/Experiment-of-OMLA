//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953;
  XNOR2_X1  g000(.A(G169gat), .B(G197gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G113gat), .B(G141gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT12), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  OR2_X1    g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n213), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT84), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT84), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n222), .B(new_n213), .C1(new_n215), .C2(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n214), .B(KEYINPUT14), .Z(new_n225));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n215), .A2(KEYINPUT86), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n219), .A2(new_n213), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT85), .B(G43gat), .Z(new_n230));
  OAI211_X1 g029(.A(new_n210), .B(new_n212), .C1(new_n230), .C2(G50gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G1gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n236), .A2(G1gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n237), .B2(new_n234), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT89), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n240), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT87), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n240), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n250), .A3(new_n232), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n224), .B2(new_n232), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n245), .A3(new_n242), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n243), .A2(new_n248), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n254), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n242), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n209), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n256), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n233), .A2(new_n240), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(new_n242), .A3(KEYINPUT89), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n233), .A3(new_n240), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n248), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n209), .A2(new_n260), .A3(new_n258), .A4(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G228gat), .ZN(new_n267));
  INV_X1    g066(.A(G233gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(G211gat), .ZN(new_n271));
  INV_X1    g070(.A(G218gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n270), .B1(KEYINPUT22), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT3), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G141gat), .B(G148gat), .Z(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT2), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n281), .A2(new_n285), .B1(new_n282), .B2(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n281), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n280), .B(new_n282), .C1(new_n289), .C2(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n269), .B1(new_n279), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI211_X1 g096(.A(KEYINPUT73), .B(KEYINPUT3), .C1(new_n287), .C2(new_n290), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT29), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n276), .B(KEYINPUT70), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n276), .B(KEYINPUT70), .Z(new_n304));
  OAI21_X1  g103(.A(new_n278), .B1(new_n296), .B2(new_n298), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT76), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n293), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G22gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(KEYINPUT75), .A3(new_n276), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT75), .B1(new_n305), .B2(new_n276), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n277), .A2(new_n278), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n291), .B1(new_n312), .B2(new_n295), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n307), .B(new_n308), .C1(new_n314), .C2(new_n269), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n276), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n269), .B1(new_n318), .B2(new_n309), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT76), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n292), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(G22gat), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n307), .B1(new_n314), .B2(new_n269), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT77), .B1(new_n325), .B2(G22gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G78gat), .B(G106gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT31), .B(G50gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n323), .A3(KEYINPUT77), .A4(new_n329), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G227gat), .A2(G233gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT64), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G183gat), .B(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n337), .B1(new_n338), .B2(new_n336), .ZN(new_n339));
  INV_X1    g138(.A(G169gat), .ZN(new_n340));
  INV_X1    g139(.A(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT65), .B(new_n337), .C1(new_n338), .C2(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n350), .B(new_n351), .C1(new_n339), .C2(new_n348), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n342), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT67), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(new_n356), .B2(new_n345), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(KEYINPUT67), .A3(new_n342), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n360), .A2(new_n361), .B1(G183gat), .B2(G190gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT27), .B(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n365), .B2(G190gat), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n364), .B(new_n367), .C1(KEYINPUT66), .C2(KEYINPUT28), .ZN(new_n368));
  NAND2_X1  g167(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G127gat), .B(G134gat), .Z(new_n373));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n374));
  INV_X1    g173(.A(G127gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n375), .A2(G134gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377));
  OAI221_X1 g176(.A(new_n373), .B1(new_n374), .B2(new_n376), .C1(KEYINPUT1), .C2(new_n377), .ZN(new_n378));
  OAI22_X1  g177(.A1(new_n377), .A2(KEYINPUT1), .B1(new_n376), .B2(new_n374), .ZN(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n372), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n382), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n355), .B2(new_n371), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n335), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G15gat), .B(G43gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n335), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n382), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n353), .A2(new_n354), .B1(new_n362), .B2(new_n370), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n384), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n392), .B1(new_n398), .B2(KEYINPUT33), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT32), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n397), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n335), .A2(KEYINPUT34), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n397), .A3(new_n334), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n404), .A2(new_n405), .B1(new_n406), .B2(KEYINPUT34), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n393), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n393), .B2(new_n402), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n333), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n287), .A2(new_n290), .A3(KEYINPUT3), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n412), .A2(new_n382), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n296), .B2(new_n298), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  INV_X1    g215(.A(new_n291), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n382), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n291), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n414), .A2(new_n415), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n382), .B(new_n291), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT5), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(new_n419), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n430), .A2(KEYINPUT5), .A3(new_n415), .A4(new_n414), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n423), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n423), .A2(new_n431), .A3(new_n428), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n434), .A2(new_n433), .A3(KEYINPUT6), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n432), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(KEYINPUT71), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n372), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n277), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n442), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n372), .A2(G226gat), .A3(G233gat), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n302), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OR4_X1    g252(.A1(KEYINPUT30), .A2(new_n445), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n449), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n444), .A3(new_n452), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n453), .B1(new_n445), .B2(new_n449), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT30), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT35), .B1(new_n411), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n423), .A2(new_n431), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT6), .B1(new_n463), .B2(new_n427), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n436), .A2(KEYINPUT78), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n423), .A2(new_n431), .A3(new_n466), .A4(new_n428), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT79), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n464), .A2(new_n465), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n432), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n459), .A2(KEYINPUT35), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n333), .A2(new_n472), .A3(new_n410), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n462), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n479), .C1(new_n408), .C2(new_n409), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n393), .A2(new_n402), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n404), .A2(new_n405), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n406), .A2(KEYINPUT34), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n393), .A2(new_n402), .A3(new_n407), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(new_n476), .A3(new_n477), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT77), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n323), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n490), .A2(new_n329), .B1(new_n315), .B2(new_n323), .ZN(new_n491));
  INV_X1    g290(.A(new_n332), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n493), .B2(new_n461), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  INV_X1    g294(.A(new_n415), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n412), .A2(new_n382), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n297), .B2(new_n299), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n498), .B2(new_n429), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n421), .B2(new_n415), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n496), .C1(new_n498), .C2(new_n429), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n427), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n495), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(new_n501), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(KEYINPUT40), .A3(new_n427), .A4(new_n503), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n465), .A2(new_n467), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n454), .A4(new_n458), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n452), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n457), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n447), .A2(new_n448), .A3(new_n302), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n277), .B1(new_n441), .B2(new_n443), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT37), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n511), .B1(new_n455), .B2(new_n444), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n457), .B2(new_n513), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n519), .B(new_n456), .C1(new_n521), .C2(new_n515), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n333), .B(new_n510), .C1(new_n472), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n494), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n266), .B1(new_n475), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT91), .B(G64gat), .ZN(new_n526));
  INV_X1    g325(.A(G57gat), .ZN(new_n527));
  OR3_X1    g326(.A1(new_n526), .A2(KEYINPUT92), .A3(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G71gat), .B(G78gat), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT9), .ZN(new_n531));
  INV_X1    g330(.A(G71gat), .ZN(new_n532));
  INV_X1    g331(.A(G78gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(G64gat), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT92), .B(new_n535), .C1(new_n526), .C2(new_n527), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n528), .A2(new_n530), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(KEYINPUT90), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n538), .B2(KEYINPUT90), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n529), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G127gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n249), .B1(new_n543), .B2(new_n542), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT93), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G155gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G183gat), .B(G211gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n550), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n557), .A2(KEYINPUT98), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT41), .ZN(new_n559));
  INV_X1    g358(.A(G232gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n268), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  INV_X1    g364(.A(G92gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(KEYINPUT95), .ZN(new_n572));
  AND2_X1   g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT94), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT7), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n568), .B(new_n572), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n569), .B1(new_n571), .B2(KEYINPUT95), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(KEYINPUT7), .A3(new_n576), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n568), .B1(new_n581), .B2(new_n572), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n567), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(new_n567), .C1(new_n579), .C2(new_n582), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT97), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n589), .A3(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n233), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n252), .A2(new_n253), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n592), .B(new_n593), .C1(new_n591), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n557), .A2(KEYINPUT98), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n595), .B2(new_n596), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n563), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n562), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n555), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n542), .A3(new_n590), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g409(.A(new_n542), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(new_n586), .A3(new_n587), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n608), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n607), .B1(new_n609), .B2(new_n612), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(KEYINPUT99), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n617), .B2(KEYINPUT99), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n615), .B2(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n606), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n525), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n439), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g431(.A1(new_n628), .A2(new_n460), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n239), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n239), .B2(new_n633), .ZN(new_n637));
  MUX2_X1   g436(.A(new_n636), .B(new_n637), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g437(.A1(new_n480), .A2(new_n487), .ZN(new_n639));
  OAI21_X1  g438(.A(G15gat), .B1(new_n628), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n410), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(G15gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n628), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n629), .A2(new_n493), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT101), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n494), .A2(new_n523), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n494), .B2(new_n523), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n475), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n648), .B1(new_n653), .B2(new_n605), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n475), .A2(new_n524), .ZN(new_n655));
  INV_X1    g454(.A(new_n605), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(KEYINPUT44), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n555), .ZN(new_n659));
  INV_X1    g458(.A(new_n626), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n259), .B2(new_n265), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n260), .A2(new_n258), .A3(new_n264), .ZN(new_n663));
  INV_X1    g462(.A(new_n209), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n209), .A2(new_n260), .A3(new_n258), .A4(new_n264), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n439), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n555), .A2(new_n605), .A3(new_n626), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n525), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(G29gat), .A3(new_n439), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT45), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(G1328gat));
  NAND2_X1  g474(.A1(new_n217), .A2(new_n218), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n669), .B2(new_n460), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n672), .A2(new_n460), .A3(new_n676), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT46), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(G1329gat));
  INV_X1    g479(.A(new_n230), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n672), .B2(new_n641), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n488), .A2(new_n230), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n669), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT47), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n686), .B(new_n682), .C1(new_n669), .C2(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1330gat));
  INV_X1    g487(.A(G50gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n672), .B2(new_n333), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n493), .A2(G50gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n669), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT48), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT48), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n694), .B(new_n690), .C1(new_n669), .C2(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n668), .A2(new_n660), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n606), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n652), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n652), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n439), .B(KEYINPUT105), .Z(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(new_n527), .ZN(G1332gat));
  AOI21_X1  g506(.A(new_n460), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1333gat));
  NOR2_X1   g512(.A1(new_n639), .A2(new_n532), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n701), .A2(new_n703), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT108), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n532), .B1(new_n704), .B2(new_n641), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n716), .B2(new_n717), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(G1334gat));
  NOR2_X1   g520(.A1(new_n704), .A2(new_n333), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n533), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n555), .A2(new_n668), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n652), .A2(KEYINPUT51), .A3(new_n656), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT110), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n472), .A2(new_n522), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n510), .B1(new_n491), .B2(new_n492), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n464), .A2(KEYINPUT74), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n436), .A3(new_n435), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n459), .B1(new_n731), .B2(new_n432), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n639), .B1(new_n333), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT103), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n494), .A2(new_n523), .A3(new_n649), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n605), .B1(new_n736), .B2(new_n475), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT51), .A4(new_n724), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n652), .A2(new_n656), .A3(new_n724), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n739), .A3(new_n742), .A4(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n565), .A3(new_n630), .A4(new_n626), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n698), .A2(new_n555), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n658), .A2(new_n630), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G85gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1336gat));
  NAND4_X1  g551(.A1(new_n654), .A2(new_n459), .A3(new_n657), .A4(new_n749), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n566), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n460), .A2(new_n660), .A3(G92gat), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(new_n743), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n753), .A2(G92gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n757), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n742), .B2(new_n725), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT52), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(G1337gat));
  NOR3_X1   g563(.A1(new_n641), .A2(new_n660), .A3(G99gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n654), .A2(new_n488), .A3(new_n657), .A4(new_n749), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G99gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(KEYINPUT113), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  INV_X1    g569(.A(new_n765), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n745), .B2(new_n746), .ZN(new_n772));
  INV_X1    g571(.A(new_n768), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n333), .A2(G106gat), .A3(new_n660), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n743), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n654), .A2(new_n493), .A3(new_n657), .A4(new_n749), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G106gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT114), .B1(new_n778), .B2(G106gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n776), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n742), .B2(new_n725), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n786), .B2(new_n780), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n613), .A2(new_n614), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n607), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n613), .A2(new_n608), .A3(new_n614), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT115), .B(new_n621), .C1(new_n615), .C2(new_n790), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n790), .A3(new_n607), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n622), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n613), .A2(new_n608), .A3(new_n614), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n615), .A3(new_n790), .ZN(new_n801));
  AOI211_X1 g600(.A(KEYINPUT54), .B(new_n608), .C1(new_n613), .C2(new_n614), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n802), .B2(new_n621), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n797), .A2(new_n796), .A3(new_n622), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n799), .B(new_n624), .C1(new_n805), .C2(KEYINPUT55), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n248), .B1(new_n262), .B2(new_n263), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n245), .B1(new_n254), .B2(new_n242), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n208), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n666), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n602), .A2(new_n604), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n788), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n811), .ZN(new_n813));
  INV_X1    g612(.A(new_n801), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n795), .B2(new_n798), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n789), .ZN(new_n816));
  INV_X1    g615(.A(new_n624), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n803), .A2(new_n804), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n794), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n813), .A2(new_n816), .A3(new_n819), .A4(KEYINPUT116), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(new_n668), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n810), .A2(new_n626), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n656), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n659), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n627), .A2(new_n667), .A3(new_n662), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n705), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n459), .A3(new_n411), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n668), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n493), .B1(new_n825), .B2(new_n826), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n630), .A2(new_n831), .A3(new_n460), .A4(new_n410), .ZN(new_n832));
  INV_X1    g631(.A(new_n266), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(G113gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n832), .B2(new_n834), .ZN(G1340gat));
  AOI21_X1  g634(.A(G120gat), .B1(new_n829), .B2(new_n626), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n626), .A2(G120gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n832), .B2(new_n837), .ZN(G1341gat));
  AOI21_X1  g637(.A(new_n375), .B1(new_n832), .B2(new_n555), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n659), .A2(G127gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n829), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT117), .ZN(G1342gat));
  NAND2_X1  g641(.A1(new_n656), .A2(new_n460), .ZN(new_n843));
  OR4_X1    g642(.A1(G134gat), .A2(new_n828), .A3(new_n411), .A4(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n832), .A2(new_n656), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G134gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(G1343gat));
  NOR3_X1   g648(.A1(new_n488), .A2(new_n439), .A3(new_n459), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n825), .A2(new_n826), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n851), .B2(new_n493), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n493), .A2(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n816), .A2(new_n819), .A3(new_n833), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n656), .B1(new_n854), .B2(new_n823), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n659), .B1(new_n821), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(new_n856), .B2(new_n826), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n850), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n266), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n639), .A2(new_n493), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n266), .A2(G141gat), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n827), .A2(new_n460), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT58), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n859), .B(new_n865), .C1(new_n864), .C2(new_n863), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n705), .B(new_n860), .C1(new_n825), .C2(new_n826), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n460), .A4(new_n862), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n668), .B(new_n850), .C1(new_n852), .C2(new_n857), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT119), .B1(new_n874), .B2(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n876), .B(new_n877), .C1(new_n871), .C2(new_n873), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n866), .B1(new_n875), .B2(new_n878), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n851), .A2(KEYINPUT57), .A3(new_n493), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n806), .A2(new_n811), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n659), .B1(new_n855), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n627), .A2(new_n266), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n333), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n880), .B1(KEYINPUT57), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n626), .A3(new_n850), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n626), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n460), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n888), .B1(new_n891), .B2(new_n626), .ZN(new_n892));
  OAI221_X1 g691(.A(new_n887), .B1(new_n858), .B2(new_n889), .C1(G148gat), .C2(new_n892), .ZN(G1345gat));
  OR3_X1    g692(.A1(new_n890), .A2(G155gat), .A3(new_n659), .ZN(new_n894));
  OAI21_X1  g693(.A(G155gat), .B1(new_n858), .B2(new_n659), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n858), .B2(new_n605), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n843), .A2(G162gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n869), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1347gat));
  AOI21_X1  g699(.A(new_n630), .B1(new_n825), .B2(new_n826), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n411), .A2(new_n460), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n340), .A3(new_n668), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n705), .A2(new_n459), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n831), .A2(new_n410), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n266), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n905), .A2(new_n341), .A3(new_n626), .ZN(new_n914));
  OAI21_X1  g713(.A(G176gat), .B1(new_n908), .B2(new_n660), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1349gat));
  OAI21_X1  g715(.A(KEYINPUT123), .B1(new_n908), .B2(new_n659), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G183gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n908), .A2(KEYINPUT123), .A3(new_n659), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n555), .A2(new_n364), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n918), .A2(new_n919), .B1(new_n903), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n908), .B2(new_n605), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n605), .A2(G190gat), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n905), .A2(KEYINPUT124), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT124), .B1(new_n905), .B2(new_n927), .ZN(new_n929));
  OAI221_X1 g728(.A(new_n926), .B1(KEYINPUT61), .B2(new_n925), .C1(new_n928), .C2(new_n929), .ZN(G1351gat));
  AND2_X1   g729(.A1(new_n907), .A2(new_n639), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n885), .A2(G197gat), .A3(new_n833), .A4(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n901), .A2(new_n459), .A3(new_n861), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n668), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n933), .A2(new_n935), .ZN(G1352gat));
  XNOR2_X1  g735(.A(KEYINPUT126), .B(G204gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n660), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT62), .Z(new_n940));
  NAND3_X1  g739(.A1(new_n885), .A2(new_n626), .A3(new_n931), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1353gat));
  NAND3_X1  g744(.A1(new_n934), .A2(new_n271), .A3(new_n555), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n885), .A2(new_n555), .A3(new_n931), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n272), .A3(new_n656), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n885), .A2(new_n656), .A3(new_n931), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n272), .ZN(G1355gat));
endmodule


