//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n219), .B(new_n221), .C1(new_n217), .C2(new_n218), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n209), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n214), .B(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT65), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n215), .A2(new_n226), .ZN(new_n227));
  AND4_X1   g026(.A1(new_n213), .A2(new_n224), .A3(new_n225), .A4(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n222), .A2(new_n209), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n231), .B(new_n212), .C1(new_n232), .C2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n212), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n242), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(new_n244), .A3(new_n238), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT68), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(KEYINPUT26), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n246), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n247), .A2(new_n248), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n243), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n230), .A2(new_n250), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n208), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT69), .B(new_n206), .C1(new_n259), .C2(KEYINPUT33), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT32), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n206), .C1(new_n259), .C2(KEYINPUT33), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(new_n261), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n206), .A2(KEYINPUT33), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n256), .A2(new_n258), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n271), .A2(new_n208), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n271), .B2(new_n208), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n262), .A2(new_n267), .A3(KEYINPUT74), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n275), .A2(new_n262), .A3(new_n267), .A4(KEYINPUT74), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT36), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  NAND2_X1  g086(.A1(new_n251), .A2(KEYINPUT77), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n230), .A2(new_n250), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT29), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n230), .A2(new_n250), .A3(new_n291), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G211gat), .A2(G218gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n298), .B2(KEYINPUT75), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n298), .A2(KEYINPUT75), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(KEYINPUT76), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n299), .A2(new_n300), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n294), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n289), .B1(new_n230), .B2(new_n250), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n291), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n251), .A2(new_n292), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n287), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT80), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n287), .C1(new_n310), .C2(new_n315), .ZN(new_n319));
  INV_X1    g118(.A(new_n287), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n288), .A2(new_n290), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n321), .A2(new_n291), .B1(new_n251), .B2(new_n292), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n320), .B(new_n309), .C1(new_n322), .C2(new_n308), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT30), .ZN(new_n324));
  INV_X1    g123(.A(new_n315), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT30), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n320), .A4(new_n309), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n317), .A2(new_n319), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G141gat), .B(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT81), .B(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(KEYINPUT82), .ZN(new_n336));
  INV_X1    g135(.A(G148gat), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n337), .A2(G141gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n336), .B(new_n333), .C1(KEYINPUT82), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G155gat), .ZN(new_n340));
  INV_X1    g139(.A(G162gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT2), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT83), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n335), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n335), .B(new_n346), .C1(new_n339), .C2(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n347), .A3(new_n255), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n344), .B2(new_n255), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n344), .A2(new_n255), .A3(new_n353), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT85), .A3(new_n354), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n351), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n344), .B(new_n255), .ZN(new_n362));
  INV_X1    g161(.A(new_n350), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n349), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n358), .A2(new_n348), .A3(new_n350), .A4(new_n354), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT0), .ZN(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  INV_X1    g171(.A(new_n366), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n360), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT6), .B(new_n372), .C1(new_n373), .C2(new_n360), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n328), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n344), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n301), .B2(new_n303), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n303), .B2(new_n301), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n382), .B2(new_n346), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n347), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n308), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G228gat), .ZN(new_n388));
  INV_X1    g187(.A(G233gat), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n383), .A2(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n308), .A3(KEYINPUT87), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n304), .A2(new_n384), .A3(new_n307), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n304), .A2(new_n307), .A3(KEYINPUT86), .A4(new_n384), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n380), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n390), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n390), .B(new_n403), .C1(new_n395), .C2(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n406), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n402), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n408), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n402), .A2(new_n404), .A3(new_n409), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n402), .B2(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n379), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n276), .B1(new_n268), .B2(KEYINPUT73), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n275), .A2(new_n262), .A3(new_n267), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(KEYINPUT36), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n282), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n376), .A2(new_n377), .A3(new_n323), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT37), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n309), .C1(new_n322), .C2(new_n308), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n287), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n325), .B2(new_n309), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT38), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n425), .A2(KEYINPUT38), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n313), .A2(new_n314), .ZN(new_n431));
  INV_X1    g230(.A(new_n308), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT89), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n322), .A2(new_n434), .A3(new_n308), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n293), .A2(new_n294), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n432), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT37), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n438), .B2(KEYINPUT37), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n430), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT91), .B(KEYINPUT38), .C1(new_n425), .C2(new_n426), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n429), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n362), .A2(new_n363), .ZN(new_n445));
  INV_X1    g244(.A(new_n348), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n357), .B2(new_n359), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT39), .B(new_n445), .C1(new_n447), .C2(new_n350), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n357), .A2(new_n359), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n348), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT39), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n363), .ZN(new_n452));
  OR2_X1    g251(.A1(KEYINPUT88), .A2(KEYINPUT40), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n448), .A2(new_n452), .A3(new_n370), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n374), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n447), .A2(new_n350), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n372), .B1(new_n456), .B2(new_n451), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n453), .B1(new_n457), .B2(new_n448), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n317), .A2(new_n319), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n324), .A2(new_n327), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n459), .A2(new_n462), .B1(new_n415), .B2(new_n411), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n415), .A2(new_n411), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n417), .A2(new_n419), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT35), .B1(new_n467), .B2(new_n379), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT92), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n379), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT35), .B1(new_n415), .B2(new_n411), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n328), .A2(KEYINPUT92), .A3(new_n378), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n280), .A4(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n421), .A2(new_n464), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G15gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(G22gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n403), .A2(G15gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT96), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n403), .A2(G15gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT96), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  AOI21_X1  g283(.A(G1gat), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n479), .B2(new_n480), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT97), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G8gat), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(KEYINPUT97), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n491), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n483), .A2(new_n484), .ZN(new_n494));
  INV_X1    g293(.A(G1gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498));
  OR2_X1    g297(.A1(G43gat), .A2(G50gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(G43gat), .A2(G50gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT94), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT94), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(G29gat), .A3(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT14), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n507), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT93), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n502), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n498), .A3(new_n500), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(new_n513), .A3(new_n511), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n519), .A2(new_n501), .A3(new_n507), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n512), .A2(G29gat), .A3(G36gat), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT14), .B1(new_n509), .B2(new_n510), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n508), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n507), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n516), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n501), .ZN(new_n528));
  INV_X1    g327(.A(new_n519), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n501), .A2(new_n507), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT95), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n492), .B(new_n497), .C1(new_n522), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(KEYINPUT17), .A3(new_n531), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n521), .B1(new_n517), .B2(new_n520), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT95), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT17), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n533), .B(new_n534), .C1(new_n538), .C2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n522), .B2(new_n532), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n497), .A2(new_n492), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n535), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n534), .A4(new_n533), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n539), .B(new_n540), .C1(new_n536), .C2(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n533), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n534), .B(KEYINPUT13), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n544), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G113gat), .B(G141gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G197gat), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT11), .B(G169gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT12), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n544), .A2(new_n549), .A3(new_n559), .A4(new_n553), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT98), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT99), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G71gat), .A3(G78gat), .ZN(new_n570));
  OR2_X1    g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G57gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G64gat), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G57gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n572), .A2(new_n580), .A3(KEYINPUT100), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT100), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n574), .A2(new_n576), .B1(new_n578), .B2(new_n567), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n567), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT101), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT101), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n589), .A3(new_n567), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n547), .B1(new_n566), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n566), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n598), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n597), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n607), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(new_n605), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n608), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n596), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n609), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n595), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(G85gat), .A3(G92gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  INV_X1    g426(.A(G85gat), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n623), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G99gat), .B(G106gat), .Z(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n539), .B2(new_n540), .ZN(new_n637));
  AND2_X1   g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n636), .A2(KEYINPUT105), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(KEYINPUT105), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n546), .A2(new_n535), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n622), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G134gat), .B(G162gat), .Z(new_n645));
  NOR2_X1   g444(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n639), .A2(new_n642), .A3(new_n622), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n647), .B(KEYINPUT106), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n643), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n592), .A2(new_n636), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n586), .A2(new_n634), .A3(new_n591), .A4(new_n635), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(new_n662), .A3(new_n658), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n586), .A2(new_n591), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n632), .B(new_n633), .Z(new_n666));
  NAND4_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .A4(KEYINPUT10), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT107), .B1(new_n658), .B2(new_n662), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n661), .B1(new_n660), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  AOI21_X1  g472(.A(KEYINPUT108), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n670), .B2(new_n673), .ZN(new_n675));
  INV_X1    g474(.A(new_n670), .ZN(new_n676));
  INV_X1    g475(.A(new_n673), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(KEYINPUT108), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n620), .A2(new_n656), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n474), .A2(new_n565), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n378), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n462), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT110), .Z(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT111), .ZN(new_n692));
  INV_X1    g491(.A(new_n681), .ZN(new_n693));
  OAI21_X1  g492(.A(G8gat), .B1(new_n693), .B2(new_n328), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(G1325gat));
  INV_X1    g494(.A(new_n420), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n281), .B2(new_n280), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n475), .B1(new_n681), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n280), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n681), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT112), .Z(G1326gat));
  INV_X1    g502(.A(new_n465), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n681), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NOR2_X1   g506(.A1(new_n474), .A2(new_n565), .ZN(new_n708));
  INV_X1    g507(.A(new_n620), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n679), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n656), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n509), .A3(new_n682), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n474), .B2(new_n656), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n464), .A2(new_n697), .A3(new_n416), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n468), .A2(new_n473), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n655), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n561), .A2(new_n562), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n378), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n714), .A2(new_n728), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n510), .A3(new_n462), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(KEYINPUT114), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n731), .A2(KEYINPUT114), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n727), .B2(new_n328), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n734), .B(new_n735), .C1(new_n732), .C2(new_n730), .ZN(G1329gat));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n698), .A3(new_n726), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n700), .A2(G43gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n708), .A2(new_n711), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n739), .B(new_n740), .C1(new_n742), .C2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n744), .B(KEYINPUT115), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n741), .A2(G43gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n737), .A3(new_n749), .A4(new_n738), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n747), .A2(new_n750), .ZN(G1330gat));
  AND4_X1   g550(.A1(G50gat), .A2(new_n723), .A3(new_n704), .A4(new_n726), .ZN(new_n752));
  AOI21_X1  g551(.A(G50gat), .B1(new_n712), .B2(new_n704), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n709), .A2(new_n724), .A3(new_n655), .ZN(new_n757));
  INV_X1    g556(.A(new_n679), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n719), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n378), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n573), .ZN(G1332gat));
  XNOR2_X1  g561(.A(new_n462), .B(KEYINPUT117), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(G1333gat));
  NOR3_X1   g567(.A1(new_n760), .A2(G71gat), .A3(new_n700), .ZN(new_n769));
  INV_X1    g568(.A(new_n760), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n698), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(G71gat), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n704), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n620), .A2(new_n724), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n656), .B1(new_n717), .B2(new_n718), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT118), .B1(new_n474), .B2(new_n656), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n780), .A2(KEYINPUT119), .A3(KEYINPUT51), .A4(new_n781), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n789), .A2(new_n628), .A3(new_n682), .A4(new_n758), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n776), .A2(new_n758), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n716), .B2(new_n722), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n378), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n763), .A2(G92gat), .A3(new_n679), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n787), .B2(new_n782), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n629), .B1(new_n792), .B2(new_n462), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n789), .A2(new_n796), .ZN(new_n801));
  INV_X1    g600(.A(new_n763), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n629), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n801), .B2(new_n804), .ZN(G1337gat));
  NOR2_X1   g604(.A1(new_n700), .A2(G99gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n758), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n793), .B2(new_n697), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1338gat));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n465), .B(new_n791), .C1(new_n716), .C2(new_n722), .ZN(new_n811));
  INV_X1    g610(.A(G106gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n465), .A2(G106gat), .A3(new_n679), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT121), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n719), .A2(new_n779), .A3(new_n655), .ZN(new_n816));
  AND4_X1   g615(.A1(KEYINPUT51), .A2(new_n781), .A3(new_n776), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n780), .B2(new_n781), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n791), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n723), .A2(new_n704), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT120), .A3(G106gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n813), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n789), .A2(new_n815), .ZN(new_n825));
  XOR2_X1   g624(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n821), .B2(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n669), .B2(new_n660), .ZN(new_n831));
  INV_X1    g630(.A(new_n660), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n663), .A2(new_n667), .A3(new_n668), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT123), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n669), .A2(new_n830), .A3(new_n660), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n677), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n677), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n831), .A2(new_n836), .A3(new_n833), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n836), .B1(new_n831), .B2(new_n833), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n670), .A2(new_n673), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n724), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n534), .B1(new_n548), .B2(new_n533), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n551), .A2(new_n552), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n558), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n675), .A2(new_n562), .A3(new_n678), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n655), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n655), .A2(new_n562), .A3(new_n853), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n840), .B1(new_n835), .B2(new_n837), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n847), .B(new_n846), .C1(new_n857), .C2(KEYINPUT55), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n709), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n757), .A2(new_n679), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n704), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n682), .A3(new_n280), .A4(new_n763), .ZN(new_n863));
  INV_X1    g662(.A(G113gat), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n863), .A2(new_n864), .A3(new_n565), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n378), .B1(new_n860), .B2(new_n861), .ZN(new_n866));
  INV_X1    g665(.A(new_n467), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n802), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n724), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n864), .B2(new_n870), .ZN(G1340gat));
  INV_X1    g670(.A(G120gat), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n863), .A2(new_n872), .A3(new_n679), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n758), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(G1341gat));
  INV_X1    g674(.A(G127gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n869), .A2(new_n876), .A3(new_n620), .ZN(new_n877));
  OAI21_X1  g676(.A(G127gat), .B1(new_n863), .B2(new_n709), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1342gat));
  OR4_X1    g678(.A1(G134gat), .A2(new_n868), .A3(new_n462), .A4(new_n656), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n863), .B2(new_n656), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  NOR3_X1   g683(.A1(new_n698), .A2(new_n378), .A3(new_n802), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n860), .A2(new_n861), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n704), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(new_n859), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n562), .A2(new_n675), .A3(new_n678), .A4(new_n853), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT98), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n724), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n562), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n849), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n895), .B2(new_n655), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n709), .ZN(new_n897));
  AOI211_X1 g696(.A(new_n888), .B(new_n465), .C1(new_n897), .C2(new_n861), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n885), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n565), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n698), .A2(new_n465), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n866), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n802), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n565), .A2(G141gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT58), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n899), .A2(new_n725), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n907), .A2(G141gat), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n903), .A2(new_n337), .A3(new_n758), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n620), .A2(new_n656), .A3(new_n565), .A4(new_n679), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n896), .B2(new_n709), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n704), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n854), .B1(new_n565), .B2(new_n858), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n859), .B1(new_n918), .B2(new_n656), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n913), .B1(new_n919), .B2(new_n620), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n888), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n465), .B1(new_n920), .B2(KEYINPUT125), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n915), .A2(new_n916), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT57), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n886), .A2(KEYINPUT57), .A3(new_n704), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n923), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n758), .B1(new_n885), .B2(KEYINPUT124), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(KEYINPUT124), .B2(new_n885), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n912), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n899), .A2(new_n679), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(new_n912), .A3(G148gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n911), .B1(new_n934), .B2(new_n936), .ZN(G1345gat));
  OAI21_X1  g736(.A(G155gat), .B1(new_n899), .B2(new_n709), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n903), .A2(new_n340), .A3(new_n620), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1346gat));
  OAI21_X1  g739(.A(G162gat), .B1(new_n899), .B2(new_n656), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n328), .A2(new_n341), .A3(new_n655), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n902), .B2(new_n942), .ZN(G1347gat));
  AOI211_X1 g742(.A(new_n682), .B(new_n763), .C1(new_n860), .C2(new_n861), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(new_n867), .ZN(new_n945));
  AOI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n724), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n462), .A2(new_n378), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n700), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n862), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n565), .A2(new_n217), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1348gat));
  INV_X1    g750(.A(new_n949), .ZN(new_n952));
  OAI21_X1  g751(.A(G176gat), .B1(new_n952), .B2(new_n679), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n945), .A2(new_n218), .A3(new_n758), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1349gat));
  OAI21_X1  g754(.A(G183gat), .B1(new_n952), .B2(new_n709), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n944), .A2(new_n867), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n620), .A2(new_n240), .A3(new_n241), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g759(.A(new_n212), .B1(new_n949), .B2(new_n655), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT61), .Z(new_n962));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n212), .A3(new_n655), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1351gat));
  NOR2_X1   g763(.A1(new_n698), .A2(new_n947), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n929), .B1(new_n926), .B2(new_n927), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT126), .B(KEYINPUT57), .C1(new_n924), .C2(new_n925), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n894), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n930), .A2(KEYINPUT127), .A3(new_n894), .A4(new_n965), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(new_n971), .A3(G197gat), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n944), .A2(new_n901), .ZN(new_n973));
  INV_X1    g772(.A(G197gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n973), .A2(new_n974), .A3(new_n724), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n972), .A2(new_n975), .ZN(G1352gat));
  INV_X1    g775(.A(G204gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n973), .A2(new_n977), .A3(new_n758), .ZN(new_n978));
  XOR2_X1   g777(.A(new_n978), .B(KEYINPUT62), .Z(new_n979));
  AND3_X1   g778(.A1(new_n930), .A2(new_n758), .A3(new_n965), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n977), .B2(new_n980), .ZN(G1353gat));
  INV_X1    g780(.A(G211gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n973), .A2(new_n982), .A3(new_n620), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n620), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n988), .A3(new_n655), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n930), .A2(new_n655), .A3(new_n965), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n988), .ZN(G1355gat));
endmodule


