//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT85), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n203), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT17), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G1gat), .B2(new_n214), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(G8gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n212), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT86), .B1(new_n211), .B2(new_n212), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT87), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n218), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(KEYINPUT18), .A3(new_n227), .A4(new_n228), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n211), .B(new_n218), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n226), .B(KEYINPUT13), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G197gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT11), .B(G169gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n231), .A2(new_n243), .A3(new_n232), .A4(new_n235), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G134gat), .B(G162gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT41), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n247), .B(new_n250), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  INV_X1    g055(.A(G92gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(KEYINPUT8), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G99gat), .B(G106gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  OAI221_X1 g060(.A(new_n261), .B1(new_n212), .B2(new_n211), .C1(new_n222), .C2(new_n223), .ZN(new_n262));
  XNOR2_X1  g061(.A(G190gat), .B(G218gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT93), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(KEYINPUT93), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n249), .B2(new_n248), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n259), .B(new_n260), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n211), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n265), .B1(new_n262), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n252), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n251), .A3(new_n270), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G78gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT9), .ZN(new_n285));
  INV_X1    g084(.A(G71gat), .ZN(new_n286));
  INV_X1    g085(.A(G78gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n282), .A2(new_n283), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n280), .B(new_n281), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n292), .A2(new_n288), .A3(new_n278), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT21), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n291), .A2(new_n294), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n218), .B1(new_n300), .B2(KEYINPUT21), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n299), .B(new_n301), .Z(new_n302));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT91), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G183gat), .B(G211gat), .Z(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT92), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n306), .B(new_n308), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n309), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n277), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n300), .A2(new_n268), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n261), .A2(new_n295), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT94), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n315), .A2(new_n317), .A3(new_n321), .A4(new_n316), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n300), .A2(KEYINPUT10), .A3(new_n268), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n314), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G176gat), .B(G204gat), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  AOI21_X1  g127(.A(new_n314), .B1(new_n315), .B2(new_n317), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT95), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n325), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n325), .B2(new_n330), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(G197gat), .A2(G204gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344));
  INV_X1    g143(.A(G211gat), .ZN(new_n345));
  INV_X1    g144(.A(G218gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n341), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n342), .B2(KEYINPUT80), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(KEYINPUT80), .B2(new_n342), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n337), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G141gat), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT74), .ZN(new_n362));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT2), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n366), .A2(new_n363), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT75), .B(G141gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n356), .B1(new_n368), .B2(new_n355), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n366), .B2(KEYINPUT2), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n365), .A2(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n371), .B2(new_n336), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n373), .A3(new_n341), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n342), .B(new_n374), .ZN(new_n375));
  OAI22_X1  g174(.A1(new_n354), .A2(new_n371), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G228gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n372), .A2(new_n375), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n350), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n371), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n382), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(G22gat), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n382), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n385), .A2(new_n380), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n388), .A2(new_n389), .B1(new_n376), .B2(new_n380), .ZN(new_n390));
  INV_X1    g189(.A(G22gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT81), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G50gat), .ZN(new_n396));
  XOR2_X1   g195(.A(G78gat), .B(G106gat), .Z(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n387), .A2(new_n392), .A3(KEYINPUT81), .A4(new_n398), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT70), .ZN(new_n405));
  INV_X1    g204(.A(G127gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(G134gat), .ZN(new_n407));
  INV_X1    g206(.A(G134gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(G127gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(G127gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(G134gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT70), .ZN(new_n413));
  INV_X1    g212(.A(G113gat), .ZN(new_n414));
  INV_X1    g213(.A(G120gat), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT1), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G113gat), .A2(G120gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n412), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n405), .A3(new_n417), .A4(new_n416), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n421), .A3(KEYINPUT76), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n421), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n422), .A2(new_n425), .B1(new_n371), .B2(new_n336), .ZN(new_n426));
  XNOR2_X1  g225(.A(G141gat), .B(G148gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n364), .B1(new_n427), .B2(KEYINPUT74), .ZN(new_n428));
  INV_X1    g227(.A(new_n362), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n367), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n369), .A2(new_n370), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT3), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n404), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT5), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n423), .A2(new_n430), .A3(new_n431), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n423), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n438), .A2(KEYINPUT78), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT78), .B1(new_n438), .B2(new_n439), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n434), .B(new_n435), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n371), .B1(new_n425), .B2(new_n422), .ZN(new_n443));
  INV_X1    g242(.A(new_n436), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n404), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n431), .A3(new_n336), .ZN(new_n446));
  INV_X1    g245(.A(new_n422), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT76), .B1(new_n419), .B2(new_n421), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n371), .A2(new_n384), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n403), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n438), .A2(new_n439), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n445), .B(KEYINPUT5), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT0), .ZN(new_n456));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n453), .A3(new_n458), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466));
  NAND3_X1  g265(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(G183gat), .B2(G190gat), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(G183gat), .ZN(new_n472));
  INV_X1    g271(.A(G190gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n474), .A3(KEYINPUT64), .A4(new_n467), .ZN(new_n475));
  INV_X1    g274(.A(G169gat), .ZN(new_n476));
  INV_X1    g275(.A(G176gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT23), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(G169gat), .B2(G176gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G169gat), .A2(G176gat), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n470), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n476), .A2(new_n477), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n487), .B2(new_n479), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(G169gat), .A3(G176gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n481), .A2(KEYINPUT65), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n488), .A2(new_n478), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT24), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n494), .B1(G183gat), .B2(G190gat), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n468), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n486), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n491), .A3(new_n490), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n480), .A2(KEYINPUT25), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G183gat), .A2(G190gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(KEYINPUT66), .B2(KEYINPUT24), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n474), .B(new_n467), .C1(new_n504), .C2(new_n495), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(KEYINPUT67), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n487), .A2(KEYINPUT26), .ZN(new_n508));
  NOR2_X1   g307(.A1(G169gat), .A2(G176gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n481), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n503), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(new_n473), .C1(new_n472), .C2(KEYINPUT27), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n515), .A2(KEYINPUT69), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT69), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n473), .B1(new_n472), .B2(KEYINPUT27), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT27), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(G183gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n519), .A2(new_n521), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n515), .A2(new_n516), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n515), .A2(KEYINPUT69), .A3(new_n516), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n513), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G226gat), .A2(G233gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n522), .B1(new_n517), .B2(new_n518), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n524), .A3(new_n528), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n512), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n478), .A2(new_n491), .A3(new_n490), .ZN(new_n536));
  AND4_X1   g335(.A1(KEYINPUT67), .A2(new_n505), .A3(new_n488), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT67), .B1(new_n502), .B2(new_n505), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(new_n485), .ZN(new_n540));
  INV_X1    g339(.A(new_n531), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(KEYINPUT29), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n375), .B(new_n532), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n507), .B2(new_n530), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n375), .A4(new_n532), .ZN(new_n548));
  INV_X1    g347(.A(new_n375), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n507), .A2(new_n530), .A3(new_n531), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  XNOR2_X1  g350(.A(G8gat), .B(G36gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G64gat), .B(G92gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n552), .B(new_n553), .Z(new_n554));
  NAND4_X1  g353(.A1(new_n544), .A2(new_n548), .A3(new_n551), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n554), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n556), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n544), .A2(new_n548), .A3(new_n551), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n548), .A3(new_n551), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n558), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n402), .B1(new_n465), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n423), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n507), .A2(new_n530), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n565), .B1(new_n507), .B2(new_n530), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G227gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT34), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT34), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n572), .B(new_n569), .C1(new_n566), .C2(new_n567), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT33), .B1(new_n568), .B2(new_n570), .ZN(new_n574));
  XNOR2_X1  g373(.A(G15gat), .B(G43gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G99gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n571), .B(new_n573), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n507), .A2(new_n530), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n423), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n507), .A2(new_n530), .A3(new_n565), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n570), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n577), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n581), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n572), .B1(new_n587), .B2(new_n569), .ZN(new_n588));
  INV_X1    g387(.A(new_n573), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n578), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n584), .B1(new_n578), .B2(new_n590), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n591), .A2(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n590), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n583), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n590), .A3(new_n584), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n551), .A2(new_n543), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT38), .B1(new_n603), .B2(KEYINPUT37), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n604), .B(new_n558), .C1(KEYINPUT37), .C2(new_n561), .ZN(new_n605));
  AND4_X1   g404(.A1(new_n464), .A2(new_n605), .A3(new_n463), .A4(new_n555), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT83), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n561), .A2(KEYINPUT37), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n558), .B1(new_n561), .B2(KEYINPUT37), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n607), .B(KEYINPUT38), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n558), .A2(KEYINPUT37), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n562), .A2(new_n611), .B1(KEYINPUT37), .B2(new_n561), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT83), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n606), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n400), .A2(new_n401), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n436), .A2(new_n437), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT4), .B1(new_n371), .B2(new_n423), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT78), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n621), .A2(new_n622), .B1(new_n433), .B2(new_n426), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT82), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n623), .A2(new_n624), .A3(new_n403), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n426), .A2(new_n433), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n440), .B2(new_n441), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT82), .B1(new_n627), .B2(new_n404), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n617), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n624), .B1(new_n623), .B2(new_n403), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(KEYINPUT82), .A3(new_n404), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n443), .A2(new_n444), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n617), .B1(new_n632), .B2(new_n403), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n629), .A2(KEYINPUT40), .A3(new_n458), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n460), .A3(new_n563), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n631), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n459), .B1(new_n637), .B2(new_n617), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT40), .B1(new_n638), .B2(new_n634), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n616), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n564), .B(new_n602), .C1(new_n615), .C2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n402), .A2(new_n591), .A3(new_n592), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT35), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n465), .A2(new_n563), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n642), .A2(KEYINPUT84), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n591), .A2(new_n592), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n616), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n563), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n463), .A2(new_n464), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT84), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT35), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n246), .B(new_n335), .C1(new_n641), .C2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n465), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n653), .A2(new_n563), .ZN(new_n657));
  INV_X1    g456(.A(G8gat), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n656), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n656), .B2(new_n661), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n653), .A2(new_n666), .A3(new_n646), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n595), .A2(new_n668), .A3(new_n601), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n595), .B2(new_n601), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n653), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n667), .B1(new_n675), .B2(new_n666), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n653), .A2(new_n402), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT99), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n641), .A2(new_n652), .ZN(new_n681));
  INV_X1    g480(.A(new_n312), .ZN(new_n682));
  INV_X1    g481(.A(new_n334), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n246), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n681), .A2(new_n277), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n206), .A3(new_n465), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n276), .A2(KEYINPUT44), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n591), .A2(new_n592), .A3(new_n599), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n593), .A2(new_n594), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n597), .B2(new_n598), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT97), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n595), .A2(new_n601), .A3(new_n668), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n606), .A2(new_n610), .A3(new_n614), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n629), .A2(new_n458), .A3(new_n634), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n699), .A2(new_n460), .A3(new_n563), .A4(new_n635), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n696), .A2(new_n616), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n694), .A2(new_n695), .A3(new_n701), .A4(new_n564), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n652), .ZN(new_n703));
  INV_X1    g502(.A(new_n564), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n635), .A2(new_n460), .A3(new_n563), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n402), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(new_n696), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n695), .B1(new_n707), .B2(new_n694), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n688), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n681), .A2(new_n277), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n684), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(new_n465), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n687), .B1(new_n714), .B2(new_n206), .ZN(G1328gat));
  NAND3_X1  g514(.A1(new_n685), .A2(new_n207), .A3(new_n563), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT101), .B(KEYINPUT46), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n713), .A2(new_n563), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n207), .ZN(G1329gat));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n685), .A2(new_n721), .A3(new_n646), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n713), .A2(new_n671), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT47), .B(new_n722), .C1(new_n723), .C2(new_n721), .ZN(new_n724));
  INV_X1    g523(.A(new_n722), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n713), .A2(new_n674), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(KEYINPUT47), .B2(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(G50gat), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n685), .A2(new_n729), .A3(new_n402), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n713), .A2(new_n402), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(KEYINPUT102), .ZN(new_n734));
  OAI21_X1  g533(.A(G50gat), .B1(new_n733), .B2(KEYINPUT102), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n733), .A2(new_n729), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n731), .B1(new_n737), .B2(new_n730), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n703), .A2(new_n708), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n313), .A2(new_n246), .A3(new_n683), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n649), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT105), .B(G57gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1332gat));
  OR2_X1    g549(.A1(new_n648), .A2(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n648), .A2(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  AND4_X1   g558(.A1(G71gat), .A2(new_n743), .A3(new_n674), .A4(new_n744), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n646), .A3(new_n744), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762));
  AOI21_X1  g561(.A(G71gat), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n743), .A2(KEYINPUT107), .A3(new_n646), .A4(new_n744), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n766), .ZN(new_n768));
  AOI211_X1 g567(.A(new_n768), .B(new_n760), .C1(new_n763), .C2(new_n764), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(G1334gat));
  NOR2_X1   g569(.A1(new_n745), .A2(new_n616), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(new_n287), .ZN(G1335gat));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n564), .B1(new_n615), .B2(new_n640), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT100), .B1(new_n774), .B2(new_n671), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n652), .A3(new_n702), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n776), .A2(new_n688), .B1(new_n710), .B2(KEYINPUT44), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n682), .A2(new_n245), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n334), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n712), .A2(KEYINPUT109), .A3(new_n780), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n649), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n778), .A2(new_n277), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n740), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT51), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n787), .A2(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(KEYINPUT110), .A3(KEYINPUT51), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n334), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n465), .A2(new_n256), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n785), .B1(new_n796), .B2(new_n797), .ZN(G1336gat));
  NOR3_X1   g597(.A1(new_n754), .A2(G92gat), .A3(new_n334), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n777), .A2(new_n754), .A3(new_n781), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(new_n801), .C1(new_n257), .C2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n782), .A2(new_n783), .A3(new_n563), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n804), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT112), .B1(new_n804), .B2(G92gat), .ZN(new_n806));
  INV_X1    g605(.A(new_n799), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n791), .B2(new_n788), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n809), .B2(new_n801), .ZN(G1337gat));
  INV_X1    g609(.A(new_n674), .ZN(new_n811));
  OAI21_X1  g610(.A(G99gat), .B1(new_n784), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n646), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n813), .A2(G99gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n796), .B2(new_n814), .ZN(G1338gat));
  NOR3_X1   g614(.A1(new_n616), .A2(new_n334), .A3(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n793), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n712), .A2(new_n402), .A3(new_n780), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  XNOR2_X1  g618(.A(KEYINPUT113), .B(G106gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n818), .B2(KEYINPUT114), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n791), .A2(new_n788), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n782), .A2(new_n783), .A3(new_n402), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n824), .A2(new_n816), .B1(new_n825), .B2(new_n820), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n823), .B2(new_n826), .ZN(G1339gat));
  NAND3_X1  g626(.A1(new_n313), .A2(new_n246), .A3(new_n334), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n314), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n322), .A2(new_n323), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n319), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n328), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n830), .A3(new_n319), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n325), .A2(new_n835), .A3(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n331), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n227), .B1(new_n224), .B2(new_n228), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n233), .A2(new_n234), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n240), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n244), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT55), .B1(new_n834), .B2(new_n836), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n276), .A2(new_n838), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n842), .A2(new_n334), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n838), .A2(new_n843), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n245), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n848), .B2(new_n277), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n829), .B1(new_n849), .B2(new_n312), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n402), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n851), .A2(new_n465), .A3(new_n646), .A4(new_n754), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n246), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n245), .ZN(new_n854));
  INV_X1    g653(.A(new_n846), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n277), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n312), .B1(new_n856), .B2(new_n844), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n828), .ZN(new_n858));
  INV_X1    g657(.A(new_n747), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n642), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n753), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n414), .A3(new_n245), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT115), .Z(G1340gat));
  NOR3_X1   g663(.A1(new_n852), .A2(new_n415), .A3(new_n334), .ZN(new_n865));
  AOI21_X1  g664(.A(G120gat), .B1(new_n861), .B2(new_n683), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  OAI21_X1  g666(.A(G127gat), .B1(new_n852), .B2(new_n312), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n861), .A2(new_n406), .A3(new_n682), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  NAND2_X1  g669(.A1(new_n277), .A2(new_n648), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n860), .A2(G134gat), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n852), .B2(new_n276), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n850), .B2(new_n747), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n858), .A2(KEYINPUT118), .A3(new_n859), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n674), .A2(new_n616), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n754), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n245), .A2(new_n357), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n694), .A2(new_n465), .A3(new_n754), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n850), .A2(new_n616), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n838), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT117), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n245), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n277), .B1(new_n895), .B2(new_n855), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n312), .B1(new_n896), .B2(new_n844), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n616), .B1(new_n897), .B2(new_n828), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n245), .B(new_n887), .C1(new_n898), .C2(new_n886), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n883), .B1(new_n899), .B2(new_n368), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n899), .B2(new_n368), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n900), .A2(new_n902), .A3(KEYINPUT58), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  AOI221_X4 g703(.A(new_n883), .B1(new_n901), .B2(new_n904), .C1(new_n899), .C2(new_n368), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n905), .ZN(G1344gat));
  OAI21_X1  g705(.A(new_n887), .B1(new_n898), .B2(new_n886), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n907), .A2(KEYINPUT59), .A3(new_n334), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT59), .B1(new_n881), .B2(new_n334), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n355), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n858), .A2(KEYINPUT57), .A3(new_n402), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT120), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n828), .B(KEYINPUT121), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n838), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n246), .B1(new_n916), .B2(KEYINPUT117), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n846), .B1(new_n917), .B2(new_n893), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n845), .B1(new_n918), .B2(new_n277), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n913), .B1(new_n919), .B2(new_n312), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n886), .B1(new_n920), .B2(new_n616), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n334), .B(new_n884), .C1(new_n912), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n908), .B(new_n910), .C1(new_n922), .C2(new_n923), .ZN(G1345gat));
  OAI21_X1  g723(.A(G155gat), .B1(new_n907), .B2(new_n312), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n312), .A2(G155gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n881), .B2(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n907), .B2(new_n276), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n871), .A2(G162gat), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n859), .A2(new_n648), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n851), .A2(new_n646), .A3(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(new_n476), .A3(new_n246), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n850), .A2(new_n465), .A3(new_n754), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(new_n642), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n245), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n476), .B2(new_n937), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n477), .A3(new_n683), .ZN(new_n939));
  OAI21_X1  g738(.A(G176gat), .B1(new_n933), .B2(new_n334), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1349gat));
  OR3_X1    g740(.A1(new_n933), .A2(KEYINPUT123), .A3(new_n312), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT123), .B1(new_n933), .B2(new_n312), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(G183gat), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n472), .A2(KEYINPUT27), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n312), .A2(new_n521), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n935), .A2(new_n642), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT122), .ZN(new_n948));
  XNOR2_X1  g747(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n944), .B2(new_n948), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n933), .B2(new_n276), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT61), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n473), .A3(new_n277), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1351gat));
  NAND3_X1  g755(.A1(new_n672), .A2(new_n673), .A3(new_n932), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n912), .B2(new_n921), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n246), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n935), .A2(new_n880), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(G197gat), .A3(new_n246), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT125), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n967), .B1(new_n959), .B2(new_n683), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n683), .A2(new_n967), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n962), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n962), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n966), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n958), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n911), .B(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n913), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n897), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT57), .B1(new_n978), .B2(new_n402), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n683), .B(new_n974), .C1(new_n976), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G204gat), .ZN(new_n981));
  INV_X1    g780(.A(new_n972), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT127), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n973), .A2(new_n983), .ZN(G1353gat));
  INV_X1    g783(.A(new_n962), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n985), .A2(new_n345), .A3(new_n682), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n682), .B(new_n974), .C1(new_n976), .C2(new_n979), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  OAI21_X1  g789(.A(G218gat), .B1(new_n960), .B2(new_n276), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n985), .A2(new_n346), .A3(new_n277), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1355gat));
endmodule


