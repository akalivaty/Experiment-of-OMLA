

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U550 ( .A1(n678), .A2(n677), .ZN(n513) );
  NOR2_X1 U551 ( .A1(n901), .A2(n613), .ZN(n622) );
  AND2_X1 U552 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U553 ( .A(n600), .B(KEYINPUT98), .ZN(n632) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n633) );
  AND2_X1 U555 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U556 ( .A1(n684), .A2(n682), .ZN(n644) );
  AND2_X1 U557 ( .A1(G160), .A2(G40), .ZN(n682) );
  AND2_X1 U558 ( .A1(n679), .A2(n513), .ZN(n680) );
  INV_X1 U559 ( .A(KEYINPUT17), .ZN(n514) );
  NAND2_X1 U560 ( .A1(n681), .A2(n680), .ZN(n722) );
  NAND2_X1 U561 ( .A1(n854), .A2(G137), .ZN(n523) );
  NOR2_X1 U562 ( .A1(G651), .A2(n567), .ZN(n768) );
  NOR2_X1 U563 ( .A1(n530), .A2(n529), .ZN(G160) );
  INV_X1 U564 ( .A(G2105), .ZN(n518) );
  AND2_X1 U565 ( .A1(n518), .A2(G2104), .ZN(n853) );
  NAND2_X1 U566 ( .A1(G102), .A2(n853), .ZN(n517) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XNOR2_X2 U568 ( .A(n515), .B(n514), .ZN(n854) );
  NAND2_X1 U569 ( .A1(G138), .A2(n854), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n517), .A2(n516), .ZN(n522) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n857) );
  NAND2_X1 U572 ( .A1(G114), .A2(n857), .ZN(n520) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n518), .ZN(n858) );
  NAND2_X1 U574 ( .A1(G126), .A2(n858), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n522), .A2(n521), .ZN(G164) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n523), .Z(n526) );
  NAND2_X1 U578 ( .A1(G101), .A2(n853), .ZN(n524) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n524), .Z(n525) );
  NAND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G113), .A2(n857), .ZN(n528) );
  NAND2_X1 U582 ( .A1(G125), .A2(n858), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U584 ( .A(G651), .ZN(n534) );
  NOR2_X1 U585 ( .A1(G543), .A2(n534), .ZN(n531) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n531), .Z(n767) );
  NAND2_X1 U587 ( .A1(G64), .A2(n767), .ZN(n533) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n567) );
  NAND2_X1 U589 ( .A1(G52), .A2(n768), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n540) );
  NOR2_X1 U591 ( .A1(n567), .A2(n534), .ZN(n772) );
  NAND2_X1 U592 ( .A1(n772), .A2(G77), .ZN(n537) );
  NOR2_X1 U593 ( .A1(G543), .A2(G651), .ZN(n535) );
  XNOR2_X1 U594 ( .A(n535), .B(KEYINPUT64), .ZN(n765) );
  NAND2_X1 U595 ( .A1(G90), .A2(n765), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U597 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U598 ( .A1(n540), .A2(n539), .ZN(G171) );
  NAND2_X1 U599 ( .A1(G89), .A2(n765), .ZN(n541) );
  XNOR2_X1 U600 ( .A(n541), .B(KEYINPUT4), .ZN(n543) );
  NAND2_X1 U601 ( .A1(G76), .A2(n772), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U603 ( .A(n544), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G63), .A2(n767), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G51), .A2(n768), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U610 ( .A1(n765), .A2(G91), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT66), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G78), .A2(n772), .ZN(n553) );
  NAND2_X1 U613 ( .A1(G53), .A2(n768), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G65), .A2(n767), .ZN(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT67), .B(n554), .ZN(n555) );
  NOR2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U619 ( .A(KEYINPUT68), .B(n559), .ZN(G299) );
  XNOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U622 ( .A1(n772), .A2(G75), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G88), .A2(n765), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G62), .A2(n767), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G50), .A2(n768), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G87), .A2(n567), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT82), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G49), .A2(n768), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n767), .A2(n571), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(G288) );
  NAND2_X1 U637 ( .A1(G61), .A2(n767), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G86), .A2(n765), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n772), .A2(G73), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n768), .A2(G48), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(G305) );
  NAND2_X1 U645 ( .A1(n772), .A2(G72), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G85), .A2(n765), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G60), .A2(n767), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G47), .A2(n768), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  OR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G290) );
  NOR2_X1 U652 ( .A1(G164), .A2(G1384), .ZN(n684) );
  NAND2_X1 U653 ( .A1(G8), .A2(n644), .ZN(n678) );
  INV_X1 U654 ( .A(G1961), .ZN(n990) );
  NAND2_X1 U655 ( .A1(n644), .A2(n990), .ZN(n588) );
  INV_X1 U656 ( .A(n644), .ZN(n596) );
  XNOR2_X1 U657 ( .A(KEYINPUT25), .B(G2078), .ZN(n929) );
  NAND2_X1 U658 ( .A1(n596), .A2(n929), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n638) );
  NOR2_X1 U660 ( .A1(G171), .A2(n638), .ZN(n594) );
  NOR2_X1 U661 ( .A1(G1966), .A2(n678), .ZN(n657) );
  NOR2_X1 U662 ( .A1(G2084), .A2(n644), .ZN(n654) );
  NOR2_X1 U663 ( .A1(n657), .A2(n654), .ZN(n589) );
  NAND2_X1 U664 ( .A1(G8), .A2(n589), .ZN(n590) );
  XNOR2_X1 U665 ( .A(KEYINPUT30), .B(n590), .ZN(n591) );
  XOR2_X1 U666 ( .A(KEYINPUT101), .B(n591), .Z(n592) );
  NOR2_X1 U667 ( .A1(G168), .A2(n592), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U669 ( .A(KEYINPUT31), .B(n595), .Z(n643) );
  INV_X1 U670 ( .A(G299), .ZN(n902) );
  NAND2_X1 U671 ( .A1(n596), .A2(G2072), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT27), .B(n597), .Z(n599) );
  NAND2_X1 U673 ( .A1(G1956), .A2(n644), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n902), .A2(n632), .ZN(n631) );
  NAND2_X1 U675 ( .A1(G56), .A2(n767), .ZN(n601) );
  XOR2_X1 U676 ( .A(KEYINPUT14), .B(n601), .Z(n607) );
  NAND2_X1 U677 ( .A1(G81), .A2(n765), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G68), .A2(n772), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT13), .B(n605), .Z(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n768), .A2(G43), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n901) );
  INV_X1 U685 ( .A(G1996), .ZN(n930) );
  OR2_X1 U686 ( .A1(n644), .A2(n930), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT26), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n644), .A2(G1341), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G66), .A2(n767), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G92), .A2(n765), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G79), .A2(n772), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G54), .A2(n768), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U697 ( .A(KEYINPUT15), .B(n620), .Z(n917) );
  NOR2_X1 U698 ( .A1(n622), .A2(n917), .ZN(n621) );
  XOR2_X1 U699 ( .A(n621), .B(KEYINPUT100), .Z(n629) );
  NAND2_X1 U700 ( .A1(n622), .A2(n917), .ZN(n627) );
  AND2_X1 U701 ( .A1(n644), .A2(G1348), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(KEYINPUT99), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n596), .A2(G2067), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n636) );
  NOR2_X1 U708 ( .A1(n902), .A2(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT29), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G171), .A2(n638), .ZN(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT97), .B(n639), .Z(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n655) );
  NAND2_X1 U715 ( .A1(n655), .A2(G286), .ZN(n652) );
  INV_X1 U716 ( .A(G8), .ZN(n650) );
  NOR2_X1 U717 ( .A1(G1971), .A2(n678), .ZN(n646) );
  NOR2_X1 U718 ( .A1(G2090), .A2(n644), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n647), .A2(G303), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(KEYINPUT102), .ZN(n649) );
  OR2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  AND2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n653), .B(KEYINPUT32), .ZN(n661) );
  NAND2_X1 U725 ( .A1(G8), .A2(n654), .ZN(n659) );
  INV_X1 U726 ( .A(n655), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n673) );
  NOR2_X1 U730 ( .A1(G1976), .A2(G288), .ZN(n903) );
  NOR2_X1 U731 ( .A1(G1971), .A2(G303), .ZN(n662) );
  NOR2_X1 U732 ( .A1(n903), .A2(n662), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n673), .A2(n663), .ZN(n664) );
  NAND2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n904) );
  NAND2_X1 U735 ( .A1(n664), .A2(n904), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n678), .A2(n665), .ZN(n666) );
  NOR2_X1 U737 ( .A1(KEYINPUT33), .A2(n666), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n903), .A2(KEYINPUT33), .ZN(n667) );
  NOR2_X1 U739 ( .A1(n667), .A2(n678), .ZN(n668) );
  NOR2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U741 ( .A(G1981), .B(G305), .Z(n920) );
  NAND2_X1 U742 ( .A1(n670), .A2(n920), .ZN(n681) );
  NOR2_X1 U743 ( .A1(G2090), .A2(G303), .ZN(n671) );
  NAND2_X1 U744 ( .A1(G8), .A2(n671), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n674), .A2(n678), .ZN(n679) );
  NOR2_X1 U747 ( .A1(G1981), .A2(G305), .ZN(n675) );
  XOR2_X1 U748 ( .A(n675), .B(KEYINPUT24), .Z(n676) );
  XNOR2_X1 U749 ( .A(KEYINPUT96), .B(n676), .ZN(n677) );
  INV_X1 U750 ( .A(n682), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n735) );
  XNOR2_X1 U752 ( .A(G2067), .B(KEYINPUT37), .ZN(n732) );
  NAND2_X1 U753 ( .A1(G104), .A2(n853), .ZN(n686) );
  NAND2_X1 U754 ( .A1(G140), .A2(n854), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U756 ( .A(KEYINPUT34), .B(n687), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n857), .A2(G116), .ZN(n688) );
  XNOR2_X1 U758 ( .A(KEYINPUT90), .B(n688), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n858), .A2(G128), .ZN(n689) );
  XOR2_X1 U760 ( .A(KEYINPUT89), .B(n689), .Z(n690) );
  NAND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U762 ( .A(n692), .B(KEYINPUT35), .Z(n693) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U764 ( .A(KEYINPUT36), .B(n695), .Z(n696) );
  XNOR2_X1 U765 ( .A(KEYINPUT91), .B(n696), .ZN(n877) );
  NOR2_X1 U766 ( .A1(n732), .A2(n877), .ZN(n968) );
  NAND2_X1 U767 ( .A1(n735), .A2(n968), .ZN(n730) );
  INV_X1 U768 ( .A(n730), .ZN(n720) );
  XNOR2_X1 U769 ( .A(G1986), .B(G290), .ZN(n908) );
  NAND2_X1 U770 ( .A1(n908), .A2(n735), .ZN(n697) );
  XNOR2_X1 U771 ( .A(n697), .B(KEYINPUT88), .ZN(n718) );
  NAND2_X1 U772 ( .A1(G107), .A2(n857), .ZN(n698) );
  XNOR2_X1 U773 ( .A(n698), .B(KEYINPUT92), .ZN(n705) );
  NAND2_X1 U774 ( .A1(G131), .A2(n854), .ZN(n700) );
  NAND2_X1 U775 ( .A1(G119), .A2(n858), .ZN(n699) );
  NAND2_X1 U776 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U777 ( .A1(G95), .A2(n853), .ZN(n701) );
  XNOR2_X1 U778 ( .A(KEYINPUT93), .B(n701), .ZN(n702) );
  NOR2_X1 U779 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U780 ( .A1(n705), .A2(n704), .ZN(n874) );
  NAND2_X1 U781 ( .A1(n874), .A2(G1991), .ZN(n715) );
  NAND2_X1 U782 ( .A1(G117), .A2(n857), .ZN(n707) );
  NAND2_X1 U783 ( .A1(G129), .A2(n858), .ZN(n706) );
  NAND2_X1 U784 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U785 ( .A1(n853), .A2(G105), .ZN(n708) );
  XOR2_X1 U786 ( .A(KEYINPUT38), .B(n708), .Z(n709) );
  NOR2_X1 U787 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U788 ( .A(n711), .B(KEYINPUT94), .ZN(n713) );
  NAND2_X1 U789 ( .A1(G141), .A2(n854), .ZN(n712) );
  NAND2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n865) );
  NAND2_X1 U791 ( .A1(n865), .A2(G1996), .ZN(n714) );
  AND2_X1 U792 ( .A1(n715), .A2(n714), .ZN(n966) );
  XNOR2_X1 U793 ( .A(KEYINPUT95), .B(n735), .ZN(n716) );
  NOR2_X1 U794 ( .A1(n966), .A2(n716), .ZN(n727) );
  INV_X1 U795 ( .A(n727), .ZN(n717) );
  NAND2_X1 U796 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n737) );
  NOR2_X1 U799 ( .A1(G1996), .A2(n865), .ZN(n723) );
  XOR2_X1 U800 ( .A(KEYINPUT103), .B(n723), .Z(n960) );
  NOR2_X1 U801 ( .A1(G1991), .A2(n874), .ZN(n970) );
  NOR2_X1 U802 ( .A1(G1986), .A2(G290), .ZN(n724) );
  XNOR2_X1 U803 ( .A(KEYINPUT104), .B(n724), .ZN(n725) );
  NOR2_X1 U804 ( .A1(n970), .A2(n725), .ZN(n726) );
  NOR2_X1 U805 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U806 ( .A1(n960), .A2(n728), .ZN(n729) );
  XNOR2_X1 U807 ( .A(KEYINPUT39), .B(n729), .ZN(n731) );
  NAND2_X1 U808 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n732), .A2(n877), .ZN(n974) );
  NAND2_X1 U810 ( .A1(n733), .A2(n974), .ZN(n734) );
  NAND2_X1 U811 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n739) );
  XOR2_X1 U813 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n738) );
  XNOR2_X1 U814 ( .A(n739), .B(n738), .ZN(G329) );
  AND2_X1 U815 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U816 ( .A(G132), .ZN(G219) );
  INV_X1 U817 ( .A(G82), .ZN(G220) );
  INV_X1 U818 ( .A(G120), .ZN(G236) );
  INV_X1 U819 ( .A(G69), .ZN(G235) );
  NAND2_X1 U820 ( .A1(G7), .A2(G661), .ZN(n740) );
  XNOR2_X1 U821 ( .A(n740), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U822 ( .A(G223), .ZN(n805) );
  NAND2_X1 U823 ( .A1(n805), .A2(G567), .ZN(n741) );
  XOR2_X1 U824 ( .A(KEYINPUT11), .B(n741), .Z(G234) );
  XOR2_X1 U825 ( .A(G860), .B(KEYINPUT70), .Z(n749) );
  NOR2_X1 U826 ( .A1(n901), .A2(n749), .ZN(n742) );
  XNOR2_X1 U827 ( .A(n742), .B(KEYINPUT71), .ZN(G153) );
  XOR2_X1 U828 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U829 ( .A1(G868), .A2(G301), .ZN(n744) );
  OR2_X1 U830 ( .A1(n917), .A2(G868), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(G284) );
  NOR2_X1 U832 ( .A1(G299), .A2(G868), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT74), .ZN(n748) );
  INV_X1 U834 ( .A(G868), .ZN(n746) );
  NOR2_X1 U835 ( .A1(n746), .A2(G286), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(G297) );
  NAND2_X1 U837 ( .A1(n749), .A2(G559), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n750), .A2(n917), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n751), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U840 ( .A1(G868), .A2(n901), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G868), .A2(n917), .ZN(n752) );
  NOR2_X1 U842 ( .A1(G559), .A2(n752), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n754), .A2(n753), .ZN(G282) );
  XOR2_X1 U844 ( .A(G2100), .B(KEYINPUT76), .Z(n764) );
  NAND2_X1 U845 ( .A1(G111), .A2(n857), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G99), .A2(n853), .ZN(n756) );
  NAND2_X1 U847 ( .A1(G135), .A2(n854), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n858), .A2(G123), .ZN(n757) );
  XOR2_X1 U850 ( .A(KEYINPUT18), .B(n757), .Z(n758) );
  NOR2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U853 ( .A(n762), .B(KEYINPUT75), .ZN(n969) );
  XNOR2_X1 U854 ( .A(G2096), .B(n969), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(G156) );
  NAND2_X1 U856 ( .A1(n765), .A2(G93), .ZN(n766) );
  XNOR2_X1 U857 ( .A(n766), .B(KEYINPUT78), .ZN(n777) );
  NAND2_X1 U858 ( .A1(G67), .A2(n767), .ZN(n770) );
  NAND2_X1 U859 ( .A1(G55), .A2(n768), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U861 ( .A(KEYINPUT80), .B(n771), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G80), .A2(n772), .ZN(n773) );
  XNOR2_X1 U863 ( .A(KEYINPUT79), .B(n773), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT81), .B(n778), .ZN(n899) );
  XOR2_X1 U867 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n779) );
  XNOR2_X1 U868 ( .A(G305), .B(n779), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n899), .B(n780), .ZN(n782) );
  XNOR2_X1 U870 ( .A(G290), .B(G299), .ZN(n781) );
  XNOR2_X1 U871 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(G303), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(G288), .ZN(n831) );
  NAND2_X1 U874 ( .A1(G559), .A2(n917), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n785), .B(n901), .ZN(n896) );
  XNOR2_X1 U876 ( .A(n831), .B(n896), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n786), .A2(G868), .ZN(n787) );
  XOR2_X1 U878 ( .A(KEYINPUT84), .B(n787), .Z(n789) );
  NOR2_X1 U879 ( .A1(n899), .A2(G868), .ZN(n788) );
  NOR2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U881 ( .A(KEYINPUT85), .B(n790), .ZN(G295) );
  NAND2_X1 U882 ( .A1(G2078), .A2(G2084), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT20), .B(n791), .Z(n792) );
  NAND2_X1 U884 ( .A1(G2090), .A2(n792), .ZN(n793) );
  XNOR2_X1 U885 ( .A(KEYINPUT21), .B(n793), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n794), .A2(G2072), .ZN(n795) );
  XNOR2_X1 U887 ( .A(KEYINPUT86), .B(n795), .ZN(G158) );
  XNOR2_X1 U888 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U889 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U890 ( .A1(G235), .A2(G236), .ZN(n796) );
  XNOR2_X1 U891 ( .A(n796), .B(KEYINPUT87), .ZN(n797) );
  NOR2_X1 U892 ( .A1(G237), .A2(n797), .ZN(n798) );
  NAND2_X1 U893 ( .A1(G108), .A2(n798), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n811), .A2(G567), .ZN(n803) );
  NOR2_X1 U895 ( .A1(G220), .A2(G219), .ZN(n799) );
  XOR2_X1 U896 ( .A(KEYINPUT22), .B(n799), .Z(n800) );
  NOR2_X1 U897 ( .A1(G218), .A2(n800), .ZN(n801) );
  NAND2_X1 U898 ( .A1(G96), .A2(n801), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n812), .A2(G2106), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n813) );
  NAND2_X1 U901 ( .A1(G661), .A2(G483), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n813), .A2(n804), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n810), .A2(G36), .ZN(G176) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n805), .ZN(G217) );
  NAND2_X1 U905 ( .A1(G15), .A2(G2), .ZN(n807) );
  INV_X1 U906 ( .A(G661), .ZN(n806) );
  NOR2_X1 U907 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U908 ( .A(n808), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n809) );
  NAND2_X1 U910 ( .A1(n810), .A2(n809), .ZN(G188) );
  NOR2_X1 U911 ( .A1(n812), .A2(n811), .ZN(G325) );
  XOR2_X1 U912 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U913 ( .A(n813), .ZN(G319) );
  XOR2_X1 U914 ( .A(G2096), .B(G2100), .Z(n815) );
  XNOR2_X1 U915 ( .A(KEYINPUT42), .B(G2678), .ZN(n814) );
  XNOR2_X1 U916 ( .A(n815), .B(n814), .ZN(n819) );
  XOR2_X1 U917 ( .A(KEYINPUT43), .B(G2090), .Z(n817) );
  XNOR2_X1 U918 ( .A(G2067), .B(G2072), .ZN(n816) );
  XNOR2_X1 U919 ( .A(n817), .B(n816), .ZN(n818) );
  XOR2_X1 U920 ( .A(n819), .B(n818), .Z(n821) );
  XNOR2_X1 U921 ( .A(G2078), .B(G2084), .ZN(n820) );
  XNOR2_X1 U922 ( .A(n821), .B(n820), .ZN(G227) );
  XOR2_X1 U923 ( .A(G1971), .B(G1961), .Z(n823) );
  XNOR2_X1 U924 ( .A(G1966), .B(G1956), .ZN(n822) );
  XNOR2_X1 U925 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U926 ( .A(n824), .B(KEYINPUT41), .Z(n826) );
  XNOR2_X1 U927 ( .A(G1986), .B(G1976), .ZN(n825) );
  XNOR2_X1 U928 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U929 ( .A(G2474), .B(G1981), .Z(n828) );
  XNOR2_X1 U930 ( .A(G1991), .B(G1996), .ZN(n827) );
  XNOR2_X1 U931 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(G229) );
  XOR2_X1 U933 ( .A(n831), .B(G286), .Z(n833) );
  XNOR2_X1 U934 ( .A(n917), .B(G171), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n834), .B(n901), .ZN(n835) );
  NOR2_X1 U937 ( .A1(G37), .A2(n835), .ZN(G397) );
  NAND2_X1 U938 ( .A1(G124), .A2(n858), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n836), .B(KEYINPUT44), .ZN(n838) );
  NAND2_X1 U940 ( .A1(n857), .A2(G112), .ZN(n837) );
  NAND2_X1 U941 ( .A1(n838), .A2(n837), .ZN(n842) );
  NAND2_X1 U942 ( .A1(G100), .A2(n853), .ZN(n840) );
  NAND2_X1 U943 ( .A1(G136), .A2(n854), .ZN(n839) );
  NAND2_X1 U944 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U945 ( .A1(n842), .A2(n841), .ZN(G162) );
  NAND2_X1 U946 ( .A1(G118), .A2(n857), .ZN(n851) );
  NAND2_X1 U947 ( .A1(n858), .A2(G130), .ZN(n843) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(n843), .ZN(n849) );
  NAND2_X1 U949 ( .A1(G106), .A2(n853), .ZN(n845) );
  NAND2_X1 U950 ( .A1(G142), .A2(n854), .ZN(n844) );
  NAND2_X1 U951 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U952 ( .A(KEYINPUT45), .B(n846), .Z(n847) );
  XNOR2_X1 U953 ( .A(KEYINPUT110), .B(n847), .ZN(n848) );
  NOR2_X1 U954 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U955 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n852), .B(G162), .ZN(n867) );
  NAND2_X1 U957 ( .A1(G103), .A2(n853), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G139), .A2(n854), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G115), .A2(n857), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G127), .A2(n858), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n953) );
  XOR2_X1 U965 ( .A(G160), .B(n953), .Z(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n876) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n869) );
  XNOR2_X1 U969 ( .A(n969), .B(KEYINPUT111), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(n870), .B(KEYINPUT113), .Z(n872) );
  XNOR2_X1 U972 ( .A(G164), .B(KEYINPUT112), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U977 ( .A1(G37), .A2(n879), .ZN(n880) );
  XNOR2_X1 U978 ( .A(KEYINPUT114), .B(n880), .ZN(G395) );
  XOR2_X1 U979 ( .A(KEYINPUT106), .B(G2446), .Z(n882) );
  XNOR2_X1 U980 ( .A(G2443), .B(G2454), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n883), .B(G2451), .Z(n885) );
  XNOR2_X1 U983 ( .A(G1348), .B(G1341), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U985 ( .A(G2435), .B(G2427), .Z(n887) );
  XNOR2_X1 U986 ( .A(G2430), .B(G2438), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(n889), .B(n888), .Z(n890) );
  NAND2_X1 U989 ( .A1(G14), .A2(n890), .ZN(n900) );
  NAND2_X1 U990 ( .A1(G319), .A2(n900), .ZN(n893) );
  NOR2_X1 U991 ( .A1(G227), .A2(G229), .ZN(n891) );
  XNOR2_X1 U992 ( .A(KEYINPUT49), .B(n891), .ZN(n892) );
  NOR2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n895) );
  NOR2_X1 U994 ( .A1(G397), .A2(G395), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(G225) );
  XNOR2_X1 U996 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U998 ( .A(G108), .ZN(G238) );
  INV_X1 U999 ( .A(G96), .ZN(G221) );
  XOR2_X1 U1000 ( .A(KEYINPUT77), .B(n896), .Z(n897) );
  NOR2_X1 U1001 ( .A1(G860), .A2(n897), .ZN(n898) );
  XNOR2_X1 U1002 ( .A(n899), .B(n898), .ZN(G145) );
  INV_X1 U1003 ( .A(n900), .ZN(G401) );
  XOR2_X1 U1004 ( .A(G16), .B(KEYINPUT56), .Z(n928) );
  XOR2_X1 U1005 ( .A(n901), .B(G1341), .Z(n916) );
  XNOR2_X1 U1006 ( .A(G1956), .B(n902), .ZN(n910) );
  INV_X1 U1007 ( .A(n903), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1009 ( .A(KEYINPUT122), .B(n906), .ZN(n907) );
  NOR2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n913) );
  XOR2_X1 U1012 ( .A(G1971), .B(G303), .Z(n911) );
  XNOR2_X1 U1013 ( .A(KEYINPUT123), .B(n911), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT124), .B(n914), .ZN(n915) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n926) );
  XOR2_X1 U1017 ( .A(G171), .B(G1961), .Z(n919) );
  XOR2_X1 U1018 ( .A(G1348), .B(n917), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G168), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(KEYINPUT57), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n952) );
  XOR2_X1 U1026 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n979) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G35), .ZN(n943) );
  XOR2_X1 U1028 ( .A(n929), .B(G27), .Z(n932) );
  XOR2_X1 U1029 ( .A(n930), .B(G32), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n938), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G25), .B(G1991), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n944) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n944), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n979), .B(n947), .ZN(n949) );
  INV_X1 U1045 ( .A(G29), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(G11), .A2(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n983) );
  XOR2_X1 U1049 ( .A(G2072), .B(n953), .Z(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(n954), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G2078), .B(G164), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(KEYINPUT119), .B(n955), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT50), .B(n958), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G2090), .B(G162), .Z(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT51), .B(n961), .Z(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n977) );
  XNOR2_X1 U1059 ( .A(G160), .B(G2084), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT116), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n972) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(KEYINPUT117), .B(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(KEYINPUT52), .B(n978), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n981), .A2(G29), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n1010) );
  XNOR2_X1 U1072 ( .A(G1986), .B(G24), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G22), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G1976), .B(G23), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT127), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(KEYINPUT58), .B(n989), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(n990), .B(G5), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n1006) );
  XOR2_X1 U1081 ( .A(G1966), .B(G21), .Z(n1004) );
  XOR2_X1 U1082 ( .A(G1956), .B(G20), .Z(n998) );
  XOR2_X1 U1083 ( .A(G1981), .B(G6), .Z(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G19), .B(G1341), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT126), .B(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT59), .B(G1348), .Z(n999) );
  XNOR2_X1 U1090 ( .A(G4), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT60), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1007), .Z(n1008) );
  NOR2_X1 U1096 ( .A1(G16), .A2(n1008), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1011), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

