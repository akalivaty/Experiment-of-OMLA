//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT90), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G122), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(KEYINPUT2), .B2(G113), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n194), .A2(KEYINPUT2), .A3(G113), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n192), .B(new_n193), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT2), .A2(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n202), .A2(new_n195), .B1(KEYINPUT2), .B2(G113), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT70), .A3(new_n192), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n203), .A2(new_n192), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n212), .B(KEYINPUT3), .C1(new_n209), .C2(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT80), .B1(new_n215), .B2(G104), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n209), .A3(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n209), .A2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n216), .A2(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n208), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n214), .A2(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT81), .A3(G101), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n214), .A2(new_n208), .A3(new_n221), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n222), .A2(KEYINPUT81), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n223), .B(new_n224), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n215), .A2(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n219), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n192), .A2(KEYINPUT5), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n233), .B(G113), .C1(KEYINPUT5), .C2(new_n235), .ZN(new_n236));
  AND4_X1   g050(.A1(new_n205), .A2(new_n227), .A3(new_n232), .A4(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n240), .B(new_n208), .C1(new_n214), .C2(new_n221), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n229), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n224), .B1(new_n245), .B2(new_n223), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n191), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n228), .A2(new_n229), .ZN(new_n248));
  INV_X1    g062(.A(new_n223), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT87), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(new_n190), .A3(new_n238), .A4(new_n230), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(new_n251), .A3(KEYINPUT6), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(new_n191), .C1(new_n239), .C2(new_n246), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT65), .A3(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n258), .A2(G146), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n258), .A2(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n271), .A3(G128), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n262), .A2(new_n270), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  INV_X1    g088(.A(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n269), .B1(new_n257), .B2(new_n259), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT0), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n263), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n277), .A2(new_n284), .B1(new_n282), .B2(new_n272), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G125), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n288), .A2(G224), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n287), .B(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n252), .A2(new_n254), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n276), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n293), .B(new_n295), .Z(new_n296));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n190), .B(KEYINPUT8), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n227), .A2(new_n232), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n205), .B2(new_n236), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n297), .B(new_n298), .C1(new_n301), .C2(new_n237), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n298), .B1(new_n301), .B2(new_n237), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT88), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n305), .B2(new_n251), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n291), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n189), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT90), .B(new_n308), .C1(new_n291), .C2(new_n306), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n291), .A2(new_n306), .A3(new_n308), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n188), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n285), .B1(new_n222), .B2(new_n207), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n228), .B2(new_n229), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n261), .A2(new_n271), .A3(new_n268), .A4(G128), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT68), .B(G128), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n268), .B1(G143), .B2(new_n256), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(new_n320), .B2(new_n277), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n319), .A2(new_n263), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n256), .A2(G143), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n269), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n317), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n227), .A2(new_n232), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n323), .A2(new_n300), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G134), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G137), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT11), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n334), .A3(G137), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n336), .ZN(new_n340));
  NAND2_X1  g154(.A1(KEYINPUT67), .A2(G137), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT11), .A2(G134), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G131), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT11), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT66), .B(G134), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(G137), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n338), .A4(new_n343), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n316), .A2(new_n330), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n288), .A2(G227), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n222), .A2(new_n207), .ZN(new_n362));
  INV_X1    g176(.A(new_n285), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n243), .B2(new_n244), .ZN(new_n365));
  INV_X1    g179(.A(new_n328), .ZN(new_n366));
  OAI22_X1  g180(.A1(new_n366), .A2(KEYINPUT10), .B1(new_n299), .B2(new_n322), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n361), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n316), .A2(new_n330), .A3(KEYINPUT83), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n351), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n353), .A2(KEYINPUT82), .A3(new_n357), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n360), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n321), .B1(new_n227), .B2(new_n232), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n351), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT12), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n353), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n356), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT84), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n372), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(G469), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n353), .A2(KEYINPUT85), .A3(new_n357), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n376), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT85), .B1(new_n353), .B2(new_n357), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT86), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n353), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n356), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n358), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n376), .A4(new_n384), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G469), .ZN(new_n395));
  INV_X1    g209(.A(G902), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(G469), .A2(G902), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n383), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT9), .B(G234), .ZN(new_n400));
  OAI21_X1  g214(.A(G221), .B1(new_n400), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(G116), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G122), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(G107), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n264), .A2(new_n266), .A3(G143), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT94), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n318), .A2(KEYINPUT94), .A3(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n258), .A2(G128), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n347), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT13), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n413), .B(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n410), .B2(new_n411), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT95), .B1(new_n419), .B2(new_n331), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT95), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n408), .A2(new_n409), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT94), .B1(new_n318), .B2(G143), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n421), .B(G134), .C1(new_n424), .C2(new_n418), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n412), .A2(KEYINPUT96), .A3(new_n347), .A4(new_n413), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n416), .A2(new_n420), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n403), .A2(KEYINPUT97), .A3(KEYINPUT14), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT97), .B1(new_n403), .B2(KEYINPUT14), .ZN(new_n430));
  OAI221_X1 g244(.A(new_n405), .B1(KEYINPUT14), .B2(new_n403), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G107), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n406), .A2(new_n215), .ZN(new_n433));
  INV_X1    g247(.A(new_n414), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n347), .B1(new_n412), .B2(new_n413), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n432), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n400), .A2(new_n437), .A3(G953), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n427), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n427), .B2(new_n436), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n396), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G237), .A2(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G214), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G143), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n445), .B(G214), .C1(new_n447), .C2(G143), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G131), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT17), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n450), .A3(new_n349), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT76), .A2(G125), .ZN(new_n456));
  INV_X1    g270(.A(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT16), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n275), .B2(G140), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n460), .A2(new_n256), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n256), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n349), .B1(new_n449), .B2(new_n450), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n455), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G113), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n209), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n458), .A2(G146), .A3(new_n459), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(KEYINPUT92), .ZN(new_n472));
  XNOR2_X1  g286(.A(G125), .B(G140), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n256), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n471), .A3(KEYINPUT92), .ZN(new_n475));
  AND4_X1   g289(.A1(KEYINPUT18), .A2(new_n449), .A3(new_n450), .A4(G131), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n449), .A2(new_n450), .B1(KEYINPUT18), .B2(G131), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n472), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n470), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n470), .B1(new_n468), .B2(new_n478), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n396), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT93), .B(new_n396), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(G475), .A3(new_n485), .ZN(new_n486));
  OAI221_X1 g300(.A(new_n396), .B1(KEYINPUT15), .B2(new_n442), .C1(new_n439), .C2(new_n440), .ZN(new_n487));
  INV_X1    g301(.A(new_n464), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT19), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n473), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n458), .A2(new_n459), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n490), .B(new_n256), .C1(new_n491), .C2(new_n489), .ZN(new_n492));
  INV_X1    g306(.A(new_n454), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n488), .B(new_n492), .C1(new_n493), .C2(new_n466), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n470), .B1(new_n478), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n468), .A2(new_n478), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n470), .ZN(new_n497));
  INV_X1    g311(.A(G475), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n396), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT20), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n478), .A2(new_n494), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n479), .B1(new_n501), .B2(new_n470), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n498), .A4(new_n396), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n444), .A2(new_n486), .A3(new_n487), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(G234), .A2(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G952), .A3(new_n288), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT21), .B(G898), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(G902), .A3(G953), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n399), .A2(new_n401), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n437), .B1(G234), .B2(new_n396), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n318), .A2(G119), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n234), .A2(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT77), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT24), .B(G110), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n318), .A2(KEYINPUT23), .A3(G119), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT23), .B1(new_n263), .B2(G119), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n234), .B2(G128), .ZN(new_n525));
  INV_X1    g339(.A(G110), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n488), .B(new_n474), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n519), .A2(new_n521), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n465), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n525), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n523), .A2(new_n525), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(G110), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n530), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n530), .B2(new_n538), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT25), .B1(new_n545), .B2(new_n396), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n530), .A2(new_n538), .ZN(new_n547));
  INV_X1    g361(.A(new_n541), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(KEYINPUT25), .A3(new_n396), .A4(new_n542), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n516), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n516), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n396), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n205), .A2(new_n206), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n351), .A2(new_n363), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n347), .A2(G137), .ZN(new_n561));
  AOI21_X1  g375(.A(G134), .B1(new_n340), .B2(new_n341), .ZN(new_n562));
  OAI21_X1  g376(.A(G131), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n350), .A2(new_n321), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT71), .B1(new_n351), .B2(new_n363), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT71), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n569), .B(new_n285), .C1(new_n345), .C2(new_n350), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(KEYINPUT30), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT72), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n575));
  NOR4_X1   g389(.A1(new_n568), .A2(new_n570), .A3(new_n572), .A4(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n567), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n560), .A2(new_n569), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n351), .A2(KEYINPUT71), .A3(new_n363), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n578), .A2(new_n559), .A3(new_n564), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n582));
  NAND2_X1  g396(.A1(new_n445), .A2(G210), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT26), .B(G101), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND4_X1  g400(.A1(new_n580), .A2(KEYINPUT74), .A3(new_n581), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n577), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n586), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n559), .B1(new_n564), .B2(new_n560), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n565), .A2(new_n558), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(KEYINPUT28), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT28), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n580), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n590), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n580), .A2(KEYINPUT74), .A3(new_n586), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n578), .A2(new_n573), .A3(new_n579), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n575), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n571), .A2(KEYINPUT72), .A3(new_n573), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n602), .B2(new_n567), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n589), .B(new_n597), .C1(new_n603), .C2(new_n581), .ZN(new_n604));
  NOR2_X1   g418(.A1(G472), .A2(G902), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n604), .A2(KEYINPUT32), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT32), .B1(new_n604), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n577), .A2(new_n590), .A3(new_n580), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n586), .B1(new_n594), .B2(new_n596), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT29), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n559), .B1(new_n571), .B2(new_n564), .ZN(new_n612));
  INV_X1    g426(.A(new_n580), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT28), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n593), .A2(KEYINPUT28), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n614), .A2(KEYINPUT29), .A3(new_n586), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n396), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n557), .B1(new_n608), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n314), .A2(new_n515), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  AND2_X1   g436(.A1(new_n399), .A2(new_n401), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n396), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT98), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n557), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n307), .A2(new_n309), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n188), .B1(new_n631), .B2(new_n313), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n439), .A2(new_n440), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n439), .A2(new_n440), .B1(KEYINPUT99), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n442), .A2(G902), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n441), .A2(new_n442), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n485), .A2(G475), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n643), .A2(new_n484), .B1(new_n500), .B2(new_n504), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n513), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n632), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n630), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NAND2_X1  g465(.A1(new_n444), .A2(new_n487), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n513), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n291), .A2(new_n306), .A3(new_n308), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n308), .B1(new_n291), .B2(new_n306), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n654), .B(new_n187), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n630), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n547), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n555), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT101), .B1(new_n552), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n549), .A2(new_n396), .A3(new_n542), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT25), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n553), .B1(new_n668), .B2(new_n550), .ZN(new_n669));
  INV_X1    g483(.A(new_n664), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n627), .A2(new_n673), .A3(new_n628), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n314), .A2(new_n515), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(KEYINPUT32), .ZN(new_n678));
  INV_X1    g492(.A(new_n598), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n581), .B1(new_n577), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n565), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n559), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n591), .B1(new_n682), .B2(new_n595), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n613), .A2(KEYINPUT28), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n586), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n587), .B1(new_n602), .B2(new_n567), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n680), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n605), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n678), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n604), .A2(KEYINPUT32), .A3(new_n605), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n619), .ZN(new_n691));
  INV_X1    g505(.A(new_n673), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n692), .A3(new_n632), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n288), .A2(G900), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(G902), .A3(new_n507), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n508), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n653), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n399), .A2(new_n401), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT103), .B(G128), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G30));
  XNOR2_X1  g518(.A(new_n698), .B(KEYINPUT39), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n623), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n312), .A2(new_n313), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT38), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n577), .A2(new_n580), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n586), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n612), .A2(new_n613), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n713), .B2(new_n590), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n625), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n606), .A2(new_n607), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n444), .A2(new_n487), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n644), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n673), .A2(new_n187), .A3(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n710), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n707), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT104), .B(G143), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G45));
  NAND3_X1  g537(.A1(new_n642), .A2(new_n645), .A3(new_n698), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n399), .A2(new_n401), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n693), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n256), .ZN(G48));
  INV_X1    g542(.A(new_n648), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n397), .A2(new_n401), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n394), .A2(new_n396), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n395), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n391), .A2(new_n376), .A3(new_n384), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n734), .A2(KEYINPUT86), .B1(new_n388), .B2(new_n356), .ZN(new_n735));
  AOI21_X1  g549(.A(G902), .B1(new_n735), .B2(new_n393), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n730), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n729), .A2(new_n620), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  INV_X1    g555(.A(new_n657), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n620), .A2(new_n742), .A3(new_n738), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  AOI21_X1  g558(.A(new_n673), .B1(new_n608), .B2(new_n619), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n514), .A3(new_n738), .A4(new_n632), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NAND3_X1  g561(.A1(new_n578), .A2(new_n564), .A3(new_n579), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n558), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n595), .B1(new_n749), .B2(new_n580), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT106), .B1(new_n750), .B2(new_n615), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n614), .A2(new_n752), .A3(new_n616), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n753), .A3(new_n590), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n680), .A2(new_n686), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n605), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n624), .A2(G472), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n552), .A2(new_n556), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n556), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT107), .B1(new_n669), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n757), .A2(new_n758), .A3(new_n512), .A4(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n718), .B(new_n187), .C1(new_n655), .C2(new_n656), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(KEYINPUT108), .A3(new_n738), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT108), .B1(new_n766), .B2(new_n738), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n404), .ZN(G24));
  NAND2_X1  g584(.A1(new_n738), .A2(new_n632), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n688), .B1(new_n754), .B2(new_n755), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n625), .B1(new_n604), .B2(new_n396), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n673), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n725), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n275), .ZN(G27));
  INV_X1    g591(.A(new_n401), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n372), .A2(new_n378), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n779), .B2(G902), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n778), .B1(new_n397), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n655), .A2(new_n188), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n312), .A2(new_n781), .A3(new_n725), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n691), .A2(new_n763), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT42), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n631), .A2(KEYINPUT90), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n656), .A2(new_n189), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n620), .A2(new_n788), .A3(new_n789), .A4(new_n781), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n349), .ZN(G33));
  NAND4_X1  g606(.A1(new_n620), .A2(new_n788), .A3(new_n700), .A4(new_n781), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT109), .B(G134), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G36));
  INV_X1    g609(.A(new_n397), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n395), .B1(new_n779), .B2(KEYINPUT45), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n380), .A2(new_n382), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n398), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n398), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n778), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n705), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n692), .B1(new_n628), .B2(new_n627), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT112), .Z(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n640), .A2(new_n641), .B1(KEYINPUT111), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n642), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n645), .B(new_n811), .C1(KEYINPUT111), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n645), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n808), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n809), .B1(new_n808), .B2(new_n818), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n788), .B(new_n806), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  OR2_X1    g636(.A1(new_n804), .A2(KEYINPUT47), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n804), .A2(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n557), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n691), .A2(new_n826), .A3(new_n724), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n788), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  INV_X1    g643(.A(new_n788), .ZN(new_n830));
  INV_X1    g644(.A(new_n730), .ZN(new_n831));
  OAI21_X1  g645(.A(G469), .B1(new_n736), .B2(KEYINPUT105), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n731), .A2(new_n732), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n830), .A2(new_n508), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n818), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT119), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n691), .A3(new_n763), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT48), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  INV_X1    g655(.A(new_n715), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n689), .A2(new_n690), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n557), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n645), .A2(new_n835), .A3(new_n642), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n763), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n846), .A2(new_n772), .A3(new_n773), .A4(new_n508), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n818), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(G952), .B(new_n288), .C1(new_n848), .C2(new_n771), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n710), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n818), .A2(new_n188), .A3(new_n738), .A4(new_n847), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n835), .A2(new_n644), .A3(new_n812), .A4(new_n844), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n837), .B2(new_n774), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n848), .A2(new_n830), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n796), .B1(new_n733), .B2(new_n737), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n778), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT117), .Z(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n825), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n858), .A2(new_n859), .A3(new_n862), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n840), .B(new_n851), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n837), .A2(new_n774), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n823), .A2(new_n824), .A3(new_n865), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n863), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n861), .A2(new_n869), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n857), .A4(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT120), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n771), .A2(new_n775), .B1(new_n693), .B2(new_n701), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n669), .A2(new_n670), .A3(new_n699), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n843), .A2(new_n632), .A3(new_n718), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n781), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n880), .A2(new_n881), .B1(new_n693), .B2(new_n726), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n878), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n878), .B2(new_n882), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n884), .A2(KEYINPUT115), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n884), .B1(KEYINPUT115), .B2(new_n885), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT114), .B1(new_n506), .B2(new_n699), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n717), .A2(new_n890), .A3(new_n644), .A4(new_n698), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n745), .A2(new_n623), .A3(new_n788), .A4(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n788), .A2(new_n774), .A3(new_n725), .A4(new_n781), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n793), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n791), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n767), .A2(new_n768), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n513), .B1(new_n646), .B2(new_n653), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n314), .A2(new_n623), .A3(new_n629), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n675), .A3(new_n746), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n620), .B(new_n738), .C1(new_n729), .C2(new_n742), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n621), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n896), .A2(new_n897), .A3(new_n901), .A4(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n888), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n769), .A2(new_n900), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n733), .A2(new_n737), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n909), .A2(new_n632), .A3(new_n831), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n673), .A2(new_n772), .A3(new_n773), .A4(new_n724), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n691), .A2(new_n632), .A3(new_n692), .ZN(new_n912));
  INV_X1    g726(.A(new_n701), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n910), .A2(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n879), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n716), .A2(new_n765), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n726), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n781), .A2(new_n916), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n918), .A3(KEYINPUT52), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n885), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n908), .A2(new_n920), .A3(new_n896), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n907), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n906), .B(KEYINPUT53), .C1(new_n887), .C2(new_n886), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT116), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n921), .A2(new_n927), .A3(new_n922), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n921), .B2(new_n922), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n925), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n877), .A2(new_n931), .B1(G952), .B2(G953), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n846), .A2(new_n188), .A3(new_n778), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT49), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n933), .B(new_n815), .C1(new_n864), .C2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT113), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n864), .A2(new_n934), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n710), .A2(new_n716), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n932), .B1(new_n936), .B2(new_n938), .ZN(G75));
  AOI21_X1  g753(.A(KEYINPUT52), .B1(new_n914), .B2(new_n918), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n884), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n922), .B1(new_n905), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT116), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n921), .A2(new_n927), .A3(new_n922), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n396), .B1(new_n945), .B2(new_n925), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G210), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n252), .A2(new_n254), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n290), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n947), .B2(new_n948), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n288), .A2(G952), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G51));
  XOR2_X1   g769(.A(new_n398), .B(KEYINPUT57), .Z(new_n956));
  INV_X1    g770(.A(new_n930), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n926), .B1(new_n945), .B2(new_n925), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(KEYINPUT121), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n394), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n799), .B(KEYINPUT122), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n946), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n954), .B1(new_n963), .B2(new_n965), .ZN(G54));
  INV_X1    g780(.A(new_n954), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n502), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n502), .B2(new_n968), .ZN(G60));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT59), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n636), .A2(new_n638), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT54), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n976), .B2(new_n930), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT123), .B1(new_n977), .B2(new_n954), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n931), .A2(new_n973), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n636), .A2(new_n638), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n977), .A2(KEYINPUT123), .A3(new_n954), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT60), .Z(new_n986));
  NAND3_X1  g800(.A1(new_n975), .A2(new_n663), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n975), .A2(new_n986), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n967), .B(new_n987), .C1(new_n988), .C2(new_n545), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT61), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G66));
  AOI21_X1  g805(.A(new_n288), .B1(new_n510), .B2(G224), .ZN(new_n992));
  INV_X1    g806(.A(new_n908), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n288), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n949), .B1(G898), .B2(new_n288), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n994), .B(new_n995), .Z(G69));
  OAI21_X1  g810(.A(new_n602), .B1(KEYINPUT30), .B2(new_n681), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n490), .B1(new_n491), .B2(new_n489), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n997), .B(new_n998), .Z(new_n999));
  NOR2_X1   g813(.A1(new_n878), .A2(new_n727), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n721), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n646), .A2(new_n653), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n620), .A2(new_n788), .A3(new_n1004), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1005), .A2(new_n706), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n828), .A2(new_n821), .A3(new_n1006), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n999), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n784), .A2(new_n765), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n804), .A2(new_n705), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AND4_X1   g827(.A1(new_n785), .A2(new_n1000), .A3(new_n790), .A4(new_n793), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n821), .A3(new_n828), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n694), .B1(new_n1015), .B2(new_n288), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1009), .B1(new_n1016), .B2(new_n999), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(G72));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  OAI21_X1  g836(.A(new_n1022), .B1(new_n1015), .B2(new_n993), .ZN(new_n1023));
  INV_X1    g837(.A(new_n609), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1020), .B1(new_n1025), .B2(new_n967), .ZN(new_n1026));
  AOI211_X1 g840(.A(KEYINPUT126), .B(new_n954), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1003), .A2(new_n1007), .A3(new_n908), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n712), .B1(new_n1028), .B2(new_n1022), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT125), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g845(.A(KEYINPUT125), .B(new_n712), .C1(new_n1028), .C2(new_n1022), .ZN(new_n1032));
  OAI22_X1  g846(.A1(new_n1026), .A2(new_n1027), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n712), .A2(new_n609), .A3(new_n1022), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n907), .B2(new_n923), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT127), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1033), .A2(new_n1036), .ZN(G57));
endmodule


