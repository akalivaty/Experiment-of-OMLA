//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT76), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  AOI21_X1  g015(.A(G128), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n200), .A2(KEYINPUT1), .A3(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n199), .A3(new_n201), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(KEYINPUT1), .A3(G146), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n208), .B(KEYINPUT78), .C1(new_n209), .C2(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G104), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(KEYINPUT77), .A3(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n215), .A2(KEYINPUT77), .A3(KEYINPUT3), .A4(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n214), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n217), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n211), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT10), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n199), .A2(new_n201), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n213), .A2(G107), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(new_n235), .B2(KEYINPUT77), .ZN(new_n236));
  INV_X1    g050(.A(new_n221), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n214), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n224), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n223), .B1(new_n220), .B2(new_n221), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n242), .B(KEYINPUT4), .C1(new_n212), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  INV_X1    g060(.A(G134), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G137), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT11), .A3(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G131), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n248), .A2(new_n250), .A3(new_n254), .A4(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n203), .B1(new_n229), .B2(new_n205), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n227), .B1(new_n258), .B2(new_n207), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n225), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n228), .A2(new_n245), .A3(new_n257), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n241), .A2(new_n244), .B1(new_n225), .B2(new_n259), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n257), .B1(new_n263), .B2(new_n228), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n196), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n207), .B(new_n208), .C1(G128), .C2(new_n209), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n225), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n225), .B2(new_n211), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n269), .B2(new_n257), .ZN(new_n270));
  INV_X1    g084(.A(new_n217), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n242), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n226), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n256), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n196), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n261), .A2(KEYINPUT79), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT79), .B1(new_n261), .B2(new_n278), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n265), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G469), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n190), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT12), .B1(new_n275), .B2(new_n256), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n266), .B(new_n257), .C1(new_n226), .C2(new_n274), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n261), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n261), .A2(new_n278), .ZN(new_n288));
  INV_X1    g102(.A(new_n264), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n196), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G469), .B1(new_n290), .B2(G902), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n192), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n194), .A2(G952), .ZN(new_n293));
  INV_X1    g107(.A(G234), .ZN(new_n294));
  INV_X1    g108(.A(G237), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n190), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT21), .B(G898), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT87), .B1(new_n200), .B2(G128), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n205), .A3(G143), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n200), .A2(G128), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n247), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT89), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n305), .A2(new_n309), .A3(new_n247), .A4(new_n306), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G122), .ZN(new_n312));
  INV_X1    g126(.A(G122), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G116), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n312), .A2(new_n314), .A3(new_n215), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n215), .B1(new_n312), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT85), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n313), .A2(G116), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n311), .A2(G122), .ZN(new_n319));
  OAI21_X1  g133(.A(G107), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT85), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n312), .A2(new_n314), .A3(new_n215), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n308), .A2(new_n310), .A3(new_n317), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT13), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n306), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n200), .A2(KEYINPUT88), .A3(KEYINPUT13), .A4(G128), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n305), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT13), .B1(new_n200), .B2(G128), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT86), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n247), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n307), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n247), .B1(new_n305), .B2(new_n306), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n322), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n312), .B1(new_n319), .B2(KEYINPUT14), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(KEYINPUT90), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT90), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n339), .B(new_n312), .C1(new_n319), .C2(KEYINPUT14), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n215), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n324), .A2(new_n332), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT91), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n317), .A2(new_n323), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n330), .B(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n305), .A2(new_n327), .A3(new_n328), .ZN(new_n347));
  OAI21_X1  g161(.A(G134), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n348), .A3(new_n310), .A4(new_n308), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT14), .B1(new_n313), .B2(G116), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT90), .B1(new_n350), .B2(new_n318), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n351), .B(new_n340), .C1(KEYINPUT14), .C2(new_n312), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G107), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n322), .C1(new_n333), .C2(new_n334), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n188), .A2(new_n357), .A3(G953), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n343), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n343), .B2(new_n356), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n190), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G478), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT15), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n366), .A2(KEYINPUT16), .A3(G140), .ZN(new_n367));
  INV_X1    g181(.A(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT16), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT72), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n372), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n198), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G125), .B(G140), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT72), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  OAI211_X1 g192(.A(G146), .B(new_n374), .C1(new_n378), .C2(new_n367), .ZN(new_n379));
  NOR2_X1   g193(.A1(G237), .A2(G953), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n381));
  AOI21_X1  g195(.A(G143), .B1(new_n380), .B2(G214), .ZN(new_n382));
  OAI21_X1  g196(.A(G131), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n295), .A2(new_n194), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n200), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n254), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT17), .B(G131), .C1(new_n381), .C2(new_n382), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n376), .A2(new_n379), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(G113), .B(G122), .Z(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT84), .B(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT18), .A2(G131), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT18), .B(G131), .C1(new_n381), .C2(new_n382), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n369), .A2(new_n370), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n369), .B2(new_n370), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n399), .A2(new_n400), .A3(G146), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n377), .A2(new_n198), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n396), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n391), .A2(new_n394), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n369), .A2(new_n370), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n377), .A2(new_n398), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT19), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(KEYINPUT19), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n198), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n383), .A2(new_n388), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n379), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n394), .B1(new_n413), .B2(new_n403), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n365), .B1(new_n404), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT20), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n365), .C1(new_n404), .C2(new_n414), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n394), .B1(new_n391), .B2(new_n403), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n190), .B1(new_n404), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n416), .A2(new_n418), .B1(G475), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n358), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n342), .A2(KEYINPUT91), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n355), .B1(new_n349), .B2(new_n354), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n343), .A2(new_n356), .A3(new_n358), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n363), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n190), .A3(new_n428), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n301), .A2(new_n364), .A3(new_n421), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n292), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n432));
  XOR2_X1   g246(.A(G116), .B(G119), .Z(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT2), .B(G113), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT2), .B(G113), .Z(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G119), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n238), .A2(new_n240), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n433), .A2(new_n434), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT5), .ZN(new_n441));
  INV_X1    g255(.A(G119), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(G116), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT80), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(new_n441), .A3(new_n442), .A4(G116), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G113), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n437), .B2(KEYINPUT5), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n440), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n244), .A2(new_n439), .B1(new_n450), .B2(new_n225), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n432), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n244), .A2(new_n439), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(new_n449), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n225), .A3(new_n438), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n432), .A3(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n234), .A2(G125), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n258), .A2(new_n366), .A3(new_n207), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G224), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G953), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n267), .A2(G125), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n366), .B1(new_n232), .B2(new_n233), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n466), .A2(new_n471), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(new_n463), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n451), .B2(new_n452), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT81), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n450), .A2(new_n478), .A3(new_n225), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n455), .A2(new_n438), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n272), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n452), .B(KEYINPUT8), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(G902), .B1(new_n476), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n468), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G210), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n468), .A2(new_n485), .A3(new_n487), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n468), .A2(new_n485), .A3(KEYINPUT82), .A4(new_n487), .ZN(new_n493));
  OAI21_X1  g307(.A(G214), .B1(G237), .B2(G902), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT83), .A4(new_n494), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n431), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n376), .A2(new_n379), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n205), .A3(G119), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n442), .A2(G128), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT24), .B(G110), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT70), .B1(new_n442), .B2(G128), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT71), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n503), .A3(new_n504), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n506), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT23), .B1(new_n205), .B2(G119), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n504), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n509), .A2(new_n512), .B1(G110), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n501), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n399), .A2(new_n400), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n511), .A2(new_n506), .ZN(new_n521));
  INV_X1    g335(.A(G110), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n514), .A2(new_n515), .A3(new_n522), .A4(new_n504), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n520), .A2(new_n198), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n379), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n501), .A2(new_n517), .B1(new_n524), .B2(new_n379), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n518), .A2(new_n525), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n190), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n529), .B1(new_n532), .B2(new_n519), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n357), .B1(G234), .B2(new_n190), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(G902), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n546), .A2(new_n547), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n232), .A2(new_n233), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n256), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT65), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT64), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n247), .B2(G137), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n249), .A2(G134), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n249), .A2(KEYINPUT64), .A3(G134), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G131), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n552), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n249), .A2(G134), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n251), .A3(new_n553), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n561), .A2(KEYINPUT65), .A3(G131), .A4(new_n557), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n559), .A2(new_n267), .A3(new_n255), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n551), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT68), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n438), .A2(new_n435), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n551), .A2(new_n563), .A3(KEYINPUT68), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n380), .A2(G210), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT27), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT26), .B(G101), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n551), .A2(new_n563), .A3(new_n568), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT66), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n567), .B1(new_n550), .B2(new_n256), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT66), .A3(new_n563), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n579), .A2(new_n581), .B1(new_n567), .B2(new_n564), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n572), .B(new_n576), .C1(new_n582), .C2(new_n571), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT30), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n551), .A2(new_n563), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n551), .B2(new_n563), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n567), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n581), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n576), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT29), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n572), .B1(new_n582), .B2(new_n571), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n576), .A2(KEYINPUT29), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n190), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G472), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n564), .A2(new_n567), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n571), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n567), .B1(new_n564), .B2(new_n565), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT28), .B1(new_n599), .B2(new_n569), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n590), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AND4_X1   g415(.A1(KEYINPUT66), .A2(new_n551), .A3(new_n563), .A4(new_n568), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT66), .B1(new_n580), .B2(new_n563), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n576), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n564), .A2(KEYINPUT30), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n551), .A2(new_n563), .A3(new_n584), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n568), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT31), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT67), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n604), .A2(new_n607), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT31), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n590), .B1(new_n579), .B2(new_n581), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n587), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n601), .A2(new_n610), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(G472), .A2(G902), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT69), .Z(new_n619));
  INV_X1    g433(.A(KEYINPUT32), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n596), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n619), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT32), .B1(new_n617), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n500), .B(new_n549), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT67), .B1(new_n615), .B2(KEYINPUT31), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n609), .B(new_n612), .C1(new_n614), .C2(new_n587), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n593), .A2(new_n590), .B1(new_n611), .B2(new_n612), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n619), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n622), .B(new_n596), .C1(new_n632), .C2(KEYINPUT32), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n500), .B1(new_n633), .B2(new_n549), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n499), .B1(new_n627), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT92), .B(G101), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  NAND2_X1  g451(.A1(new_n617), .A2(new_n624), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n630), .B2(new_n631), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n284), .A2(new_n291), .ZN(new_n642));
  INV_X1    g456(.A(new_n192), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT25), .B1(new_n544), .B2(new_n190), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n539), .B(G902), .C1(new_n543), .C2(new_n536), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n547), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n544), .A2(new_n548), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n641), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n425), .B2(new_n426), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT95), .B1(new_n651), .B2(G478), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n361), .A2(new_n653), .A3(new_n362), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n427), .B1(KEYINPUT94), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n425), .A2(new_n426), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n657), .A2(G478), .A3(new_n190), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n421), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT93), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n489), .A2(new_n665), .A3(new_n491), .ZN(new_n666));
  INV_X1    g480(.A(new_n494), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n487), .B1(new_n468), .B2(new_n485), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(KEYINPUT93), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n666), .A2(new_n301), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n664), .A2(KEYINPUT96), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT96), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n486), .A2(KEYINPUT93), .A3(new_n488), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n491), .A2(new_n665), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n494), .B(new_n673), .C1(new_n674), .C2(new_n668), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n300), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n421), .B1(new_n655), .B2(new_n661), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n650), .B1(new_n671), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT34), .B(G104), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  INV_X1    g495(.A(new_n675), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n364), .A2(new_n429), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n420), .A2(G475), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT97), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n416), .A2(new_n418), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n301), .A2(new_n682), .A3(new_n683), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n650), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT35), .B(G107), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  NOR2_X1   g508(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n535), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n548), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT98), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n699), .A3(new_n548), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n546), .B2(new_n547), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n641), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n499), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT37), .B(G110), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G12));
  NAND2_X1  g520(.A1(new_n638), .A2(new_n620), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n588), .A2(new_n597), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n600), .B1(new_n708), .B2(KEYINPUT28), .ZN(new_n709));
  INV_X1    g523(.A(new_n594), .ZN(new_n710));
  AOI21_X1  g524(.A(G902), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n583), .A2(new_n591), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n713), .A2(G472), .B1(new_n617), .B2(new_n621), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n702), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n683), .ZN(new_n716));
  INV_X1    g530(.A(G900), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n297), .B1(new_n298), .B2(new_n717), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n716), .A2(new_n687), .A3(new_n689), .A4(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n292), .A3(new_n719), .A4(new_n682), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  NAND2_X1  g535(.A1(new_n492), .A2(new_n493), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT38), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n589), .A2(new_n576), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n725), .B(new_n190), .C1(new_n576), .C2(new_n708), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n617), .A2(new_n621), .B1(G472), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n707), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n700), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n699), .B1(new_n696), .B2(new_n548), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n647), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n421), .B1(new_n364), .B2(new_n429), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n734), .A3(new_n667), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n724), .A2(new_n728), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT99), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n718), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n292), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(KEYINPUT40), .Z(new_n742));
  NAND2_X1  g556(.A1(new_n736), .A2(new_n737), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT101), .B(G143), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G45));
  AOI211_X1 g560(.A(new_n421), .B(new_n718), .C1(new_n655), .C2(new_n661), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n715), .A2(new_n292), .A3(new_n682), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  AOI21_X1  g563(.A(new_n649), .B1(new_n714), .B2(new_n707), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n282), .A2(new_n190), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT102), .A3(new_n284), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT102), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n754), .A3(G469), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n191), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n750), .B(new_n756), .C1(new_n671), .C2(new_n678), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NAND3_X1  g573(.A1(new_n691), .A2(new_n750), .A3(new_n756), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  AOI211_X1 g575(.A(new_n191), .B(new_n675), .C1(new_n753), .C2(new_n755), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n430), .A3(new_n715), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  INV_X1    g578(.A(KEYINPUT104), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n639), .B2(new_n640), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n617), .A2(new_n190), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT104), .A3(G472), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n601), .A2(new_n608), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT103), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT103), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n601), .A2(new_n771), .A3(new_n608), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n772), .A3(new_n613), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n766), .A2(new_n768), .B1(new_n624), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n649), .A2(KEYINPUT105), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n647), .A2(new_n776), .A3(new_n648), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n734), .A2(new_n300), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n762), .A2(new_n774), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  NAND3_X1  g595(.A1(new_n756), .A2(new_n682), .A3(new_n747), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n773), .A2(new_n624), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT104), .B1(new_n767), .B2(G472), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n765), .B(new_n640), .C1(new_n617), .C2(new_n190), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n783), .B(new_n732), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT106), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n766), .A2(new_n768), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n732), .A4(new_n783), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n782), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT107), .B(G125), .Z(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G27));
  AOI21_X1  g607(.A(new_n191), .B1(new_n284), .B2(new_n291), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n667), .B1(new_n492), .B2(new_n493), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n750), .A2(new_n747), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n794), .ZN(new_n799));
  INV_X1    g613(.A(new_n718), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n662), .A2(new_n663), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n775), .A2(new_n777), .B1(new_n707), .B2(new_n714), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT42), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  NAND4_X1  g620(.A1(new_n633), .A2(new_n549), .A3(new_n794), .A4(new_n795), .ZN(new_n807));
  INV_X1    g621(.A(new_n719), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n247), .ZN(G36));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n662), .B2(new_n421), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n662), .A2(new_n421), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(KEYINPUT43), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n641), .A2(new_n732), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT108), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT108), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n812), .B(new_n814), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT44), .ZN(new_n819));
  INV_X1    g633(.A(new_n284), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n290), .A2(KEYINPUT45), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n290), .A2(KEYINPUT45), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(G469), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(G469), .A2(G902), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT46), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n191), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(new_n740), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n795), .B(KEYINPUT109), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n819), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n818), .A2(KEYINPUT44), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(new_n249), .ZN(G39));
  AND2_X1   g650(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n837));
  NOR2_X1   g651(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n829), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n191), .B(new_n837), .C1(new_n827), .C2(new_n828), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n795), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n843), .A2(new_n633), .A3(new_n549), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n747), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G140), .ZN(G42));
  NAND2_X1  g660(.A1(new_n753), .A2(new_n755), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT49), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n728), .A2(new_n813), .A3(new_n667), .A4(new_n192), .ZN(new_n849));
  INV_X1    g663(.A(new_n724), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n778), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n799), .A2(new_n801), .A3(new_n797), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n803), .A2(new_n853), .B1(new_n796), .B2(new_n797), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n747), .A2(new_n794), .A3(new_n795), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n787), .B2(new_n790), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n633), .A2(new_n292), .A3(new_n732), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n795), .A2(new_n690), .A3(new_n716), .A4(new_n800), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n807), .A2(new_n808), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n854), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n757), .A2(new_n780), .A3(new_n760), .A4(new_n763), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT111), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n549), .B1(new_n623), .B2(new_n625), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT75), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n626), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n499), .B1(new_n865), .B2(new_n703), .ZN(new_n866));
  MUX2_X1   g680(.A(new_n683), .B(new_n662), .S(new_n663), .Z(new_n867));
  NAND2_X1  g681(.A1(new_n497), .A2(new_n498), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n650), .A2(new_n867), .A3(new_n868), .A4(new_n301), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n862), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n635), .A2(new_n869), .A3(new_n862), .A4(new_n704), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n860), .B(new_n861), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n787), .A2(new_n790), .ZN(new_n874));
  INV_X1    g688(.A(new_n782), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n733), .A2(new_n666), .A3(new_n669), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n707), .B2(new_n727), .ZN(new_n878));
  INV_X1    g692(.A(new_n191), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n642), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n647), .A2(new_n731), .A3(new_n800), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT113), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n702), .A2(new_n794), .A3(new_n883), .A4(new_n800), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n720), .A2(new_n748), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n876), .A2(new_n886), .A3(KEYINPUT52), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n720), .A2(new_n748), .A3(new_n885), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n791), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n852), .B1(new_n873), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  INV_X1    g708(.A(new_n859), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n805), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n757), .A2(new_n780), .A3(new_n760), .A4(new_n763), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n856), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n635), .A2(new_n869), .A3(new_n704), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT111), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n871), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n891), .A3(KEYINPUT53), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT115), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n893), .A2(new_n905), .A3(new_n894), .A4(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n870), .A2(new_n872), .ZN(new_n908));
  INV_X1    g722(.A(new_n856), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n859), .B1(new_n798), .B2(new_n804), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n861), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT112), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n898), .A2(new_n913), .A3(new_n901), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n914), .A3(new_n891), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n852), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n908), .A2(new_n911), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT114), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n902), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n894), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT116), .B1(new_n907), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n774), .A2(new_n778), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n814), .A2(new_n296), .A3(new_n812), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n762), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n293), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT117), .B1(new_n756), .B2(new_n795), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n296), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n756), .A2(KEYINPUT117), .A3(new_n795), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n728), .A2(new_n649), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n927), .B1(new_n932), .B2(new_n677), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n814), .A2(new_n812), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n934), .A3(new_n930), .ZN(new_n935));
  INV_X1    g749(.A(new_n803), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(KEYINPUT48), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n935), .A2(KEYINPUT48), .A3(new_n936), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n925), .A2(new_n832), .A3(new_n924), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n643), .B1(new_n753), .B2(new_n755), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n842), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n847), .A2(new_n879), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n724), .A2(new_n944), .A3(new_n494), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n924), .A3(new_n925), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT50), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n945), .A2(KEYINPUT50), .A3(new_n924), .A4(new_n925), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n929), .A2(new_n874), .A3(new_n934), .A4(new_n930), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n943), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT51), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n655), .A2(new_n661), .A3(new_n421), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n929), .A2(new_n930), .A3(new_n931), .A4(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n952), .A2(new_n953), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n943), .A2(new_n950), .A3(new_n960), .A4(new_n951), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT51), .B1(new_n962), .B2(new_n958), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n940), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT119), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n902), .B(KEYINPUT114), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n892), .B1(new_n873), .B2(KEYINPUT112), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT53), .B1(new_n968), .B2(new_n914), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT54), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT116), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(new_n971), .A3(new_n904), .A4(new_n906), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n923), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(G952), .A2(G953), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n851), .B1(new_n973), .B2(new_n974), .ZN(G75));
  AOI21_X1  g789(.A(new_n190), .B1(new_n893), .B2(new_n902), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT56), .B1(new_n976), .B2(G210), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n460), .A2(new_n461), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n467), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT55), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n194), .A2(G952), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n977), .B2(new_n980), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n981), .A2(new_n984), .A3(KEYINPUT120), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT120), .B1(new_n981), .B2(new_n984), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G51));
  NAND2_X1  g801(.A1(new_n893), .A2(new_n902), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT54), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n903), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n824), .B(KEYINPUT121), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT57), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n282), .B(KEYINPUT122), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n976), .A2(G469), .A3(new_n822), .A4(new_n821), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n982), .B1(new_n995), .B2(new_n996), .ZN(G54));
  AND3_X1   g811(.A1(new_n976), .A2(KEYINPUT58), .A3(G475), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n404), .A2(new_n414), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n983), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n999), .B2(new_n998), .ZN(G60));
  NAND2_X1  g815(.A1(G478), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT59), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n990), .A2(new_n660), .A3(new_n657), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n983), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n923), .A2(new_n972), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1004), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n657), .A2(new_n660), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(G63));
  XNOR2_X1  g824(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G217), .A2(G902), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n893), .B2(new_n902), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n983), .B1(new_n1014), .B2(new_n544), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n696), .B2(new_n1014), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g831(.A(G953), .B1(new_n299), .B2(new_n465), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n908), .A2(new_n897), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n978), .B1(G898), .B2(new_n194), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G69));
  NOR2_X1   g836(.A1(new_n585), .A2(new_n586), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n409), .A2(new_n410), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1023), .B(new_n1024), .Z(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(G900), .B2(G953), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n720), .A2(new_n748), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n876), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n830), .A2(new_n682), .A3(new_n733), .A4(new_n803), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n854), .A2(new_n809), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n845), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n835), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1027), .B1(new_n1034), .B2(new_n194), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1025), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n744), .A2(new_n1029), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n744), .A2(KEYINPUT62), .A3(new_n1029), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n835), .ZN(new_n1043));
  OR2_X1    g857(.A1(new_n867), .A2(KEYINPUT124), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n867), .A2(KEYINPUT124), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n843), .A2(new_n741), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1044), .A2(new_n865), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n1042), .A2(new_n1043), .A3(new_n845), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1037), .B1(new_n1048), .B2(new_n194), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1036), .B1(new_n1049), .B2(KEYINPUT125), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT126), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1049), .A2(KEYINPUT125), .ZN(new_n1054));
  NAND4_X1  g868(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1056));
  OR2_X1    g870(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1054), .ZN(new_n1058));
  OAI211_X1 g872(.A(new_n1056), .B(new_n1057), .C1(new_n1058), .C2(new_n1050), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n1055), .A2(new_n1059), .ZN(G72));
  INV_X1    g874(.A(new_n725), .ZN(new_n1061));
  NOR2_X1   g875(.A1(new_n589), .A2(new_n576), .ZN(new_n1062));
  NAND2_X1  g876(.A1(G472), .A2(G902), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1063), .B(KEYINPUT63), .Z(new_n1064));
  INV_X1    g878(.A(new_n1064), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1066), .B1(new_n967), .B2(new_n969), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1065), .B1(new_n1034), .B2(new_n1019), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n1067), .B(new_n983), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g884(.A(new_n1019), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n1064), .B1(new_n1048), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1072), .A2(new_n1061), .ZN(new_n1073));
  OR2_X1    g887(.A1(new_n1073), .A2(KEYINPUT127), .ZN(new_n1074));
  NAND2_X1  g888(.A1(new_n1073), .A2(KEYINPUT127), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(G57));
endmodule


