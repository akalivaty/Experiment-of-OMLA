//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n441, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n461), .A2(new_n463), .A3(G101), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT3), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n477), .A3(G2104), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n473), .A2(G137), .A3(new_n464), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n470), .B1(KEYINPUT70), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(new_n463), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n460), .B1(KEYINPUT69), .B2(new_n476), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(KEYINPUT3), .B1(new_n482), .B2(new_n475), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n483), .A2(new_n484), .A3(G137), .A4(new_n464), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n483), .A2(new_n464), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  OR2_X1    g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n490), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  NAND4_X1  g072(.A1(new_n473), .A2(G138), .A3(new_n464), .A4(new_n478), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n464), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n468), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n478), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n503), .A2(KEYINPUT72), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(new_n502), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n511), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n512), .B2(new_n507), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(G164));
  NOR2_X1   g089(.A1(KEYINPUT73), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n516), .A2(KEYINPUT73), .A3(KEYINPUT5), .A4(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(G543), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n524), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(new_n529), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G51), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n521), .A2(G89), .A3(new_n525), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(KEYINPUT75), .A3(new_n539), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n523), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n526), .A2(new_n547), .B1(new_n548), .B2(new_n529), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT76), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n523), .B1(new_n551), .B2(KEYINPUT76), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n526), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G81), .B1(G43), .B2(new_n533), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  AOI22_X1  g139(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n523), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n555), .A2(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(KEYINPUT77), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n572));
  MUX2_X1   g147(.A(new_n571), .B(new_n570), .S(new_n572), .Z(new_n573));
  NAND3_X1  g148(.A1(new_n566), .A2(new_n567), .A3(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n542), .A2(new_n543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(new_n535), .ZN(G286));
  NAND2_X1  g152(.A1(new_n555), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n533), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT79), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n521), .B2(G61), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n523), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n526), .A2(new_n587), .B1(new_n588), .B2(new_n529), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n555), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n523), .B2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G171), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n555), .A2(new_n598), .A3(G92), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT81), .B1(new_n526), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n519), .A2(new_n520), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n604), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n597), .B1(new_n612), .B2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(KEYINPUT80), .B2(new_n596), .ZN(G284));
  OAI21_X1  g190(.A(new_n614), .B1(KEYINPUT80), .B2(new_n596), .ZN(G321));
  NAND2_X1  g191(.A1(G299), .A2(new_n595), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n595), .B2(G168), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n595), .B2(G168), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n612), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g200(.A1(new_n481), .A2(G2105), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n468), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(KEYINPUT84), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n632), .A2(KEYINPUT84), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n637), .B1(new_n491), .B2(new_n638), .C1(new_n639), .C2(new_n488), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  OAI211_X1 g216(.A(new_n635), .B(new_n641), .C1(new_n633), .C2(new_n631), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2443), .Z(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT85), .Z(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n669), .A2(KEYINPUT17), .A3(new_n666), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n669), .B2(KEYINPUT17), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n670), .A2(new_n671), .A3(new_n665), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n677), .A3(new_n680), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n685), .C1(new_n677), .C2(new_n684), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n688), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G23), .ZN(new_n706));
  INV_X1    g281(.A(G288), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G290), .ZN(new_n716));
  OAI21_X1  g291(.A(G16), .B1(new_n716), .B2(KEYINPUT88), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(KEYINPUT88), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n697), .A2(G24), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT87), .ZN(new_n720));
  OAI21_X1  g295(.A(G1986), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n718), .A2(G1986), .A3(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n489), .A2(G119), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n492), .A2(G131), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n464), .A2(G107), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G25), .B(new_n727), .S(G29), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n714), .A2(new_n715), .A3(new_n721), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT36), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  AOI22_X1  g312(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G139), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n737), .B1(new_n738), .B2(new_n464), .C1(new_n491), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT95), .B(G2072), .Z(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n640), .A2(new_n734), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT30), .B(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n746), .A2(new_n734), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n697), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT98), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT23), .ZN(new_n753));
  INV_X1    g328(.A(G299), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n697), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n734), .B1(KEYINPUT24), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(KEYINPUT24), .B2(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n486), .B2(G29), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n750), .B(new_n756), .C1(new_n757), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n734), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n734), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT29), .Z(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n697), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n697), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(G2090), .B1(G1966), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n492), .A2(G141), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n489), .A2(G129), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT26), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n626), .A2(G105), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n771), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n770), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G171), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G5), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AND4_X1   g362(.A1(new_n769), .A2(new_n782), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n734), .A2(G27), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G164), .B2(new_n734), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT97), .B(G2078), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n761), .A2(new_n768), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n697), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n558), .B2(new_n697), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NOR2_X1   g371(.A1(new_n760), .A2(new_n757), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT96), .Z(new_n798));
  OAI211_X1 g373(.A(new_n796), .B(new_n798), .C1(new_n791), .C2(new_n790), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n697), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n612), .B2(new_n697), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT91), .B(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G2090), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n734), .A2(G26), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT93), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT28), .ZN(new_n807));
  OR2_X1    g382(.A1(G104), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n809));
  INV_X1    g384(.A(G140), .ZN(new_n810));
  INV_X1    g385(.A(G128), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n809), .B1(new_n491), .B2(new_n810), .C1(new_n811), .C2(new_n488), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT92), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(G29), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT94), .B(G2067), .Z(new_n815));
  AOI22_X1  g390(.A1(new_n764), .A2(new_n804), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n793), .A2(new_n799), .A3(new_n803), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n733), .A2(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  AOI22_X1  g395(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n523), .B1(new_n821), .B2(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n607), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n526), .A2(new_n829), .B1(new_n830), .B2(new_n529), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n831), .B1(new_n822), .B2(new_n827), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT100), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n557), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n558), .A2(new_n836), .A3(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n612), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n833), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  NAND2_X1  g424(.A1(new_n489), .A2(G130), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n492), .A2(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n464), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT101), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n727), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n629), .Z(new_n857));
  NOR2_X1   g432(.A1(new_n512), .A2(new_n507), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n778), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n813), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n740), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n857), .B(new_n861), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n496), .B(new_n640), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n486), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n864), .B1(new_n868), .B2(new_n861), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n861), .B2(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g447(.A1(new_n605), .A2(new_n610), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT10), .B1(new_n599), .B2(new_n601), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n754), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n604), .A2(G299), .A3(new_n605), .A4(new_n610), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT103), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n611), .A2(new_n879), .A3(new_n754), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(new_n876), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n877), .A2(new_n886), .A3(new_n878), .A4(new_n880), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n840), .B(new_n622), .ZN(new_n889));
  MUX2_X1   g464(.A(new_n888), .B(new_n883), .S(new_n889), .Z(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(G303), .B(G305), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n707), .B(G290), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n891), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n892), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(G868), .B2(new_n836), .ZN(G295));
  OAI21_X1  g476(.A(new_n900), .B1(G868), .B2(new_n836), .ZN(G331));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n905));
  NAND2_X1  g480(.A1(G301), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n546), .A2(new_n549), .A3(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(G286), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(G171), .A2(KEYINPUT106), .ZN(new_n910));
  OAI21_X1  g485(.A(G168), .B1(new_n910), .B2(new_n907), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n838), .A2(new_n839), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n838), .A2(new_n839), .B1(new_n909), .B2(new_n911), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(new_n884), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n912), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n915), .B1(new_n888), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n895), .B(new_n918), .C1(new_n921), .C2(new_n917), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(new_n866), .ZN(new_n923));
  INV_X1    g498(.A(new_n895), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n888), .A2(new_n920), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n917), .B1(new_n925), .B2(new_n916), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n915), .A2(KEYINPUT107), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n904), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n877), .A2(KEYINPUT41), .A3(new_n880), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n884), .A2(new_n878), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n930), .B(new_n931), .C1(new_n913), .C2(new_n914), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n920), .A2(new_n934), .A3(new_n930), .A4(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n935), .A3(new_n916), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n924), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n922), .A2(new_n937), .A3(new_n866), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n903), .B1(new_n929), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n903), .B1(new_n938), .B2(KEYINPUT43), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n928), .A2(new_n922), .A3(new_n904), .A4(new_n866), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n941), .A2(KEYINPUT109), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT109), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n940), .B(KEYINPUT110), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G397));
  INV_X1    g524(.A(G2067), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n813), .B(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n778), .B(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n727), .B(new_n729), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n480), .A2(new_n957), .A3(G40), .A4(new_n485), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n959));
  AND2_X1   g534(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n960));
  NOR2_X1   g535(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n961));
  OAI21_X1  g536(.A(G125), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n466), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n963), .A2(G2105), .B1(new_n626), .B2(G101), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n959), .A2(new_n964), .A3(new_n485), .A4(G40), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n958), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n512), .B2(new_n507), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n956), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  AND2_X1   g551(.A1(G290), .A2(G1986), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n586), .A2(new_n590), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(G1981), .B1(new_n585), .B2(new_n589), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT49), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT49), .B1(new_n982), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n503), .B2(new_n508), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n967), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(G8), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n707), .A2(G1976), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n988), .A2(G8), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n988), .A2(G8), .A3(new_n990), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n989), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(G303), .A2(G8), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n998));
  OR2_X1    g573(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n998), .B(new_n999), .Z(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n958), .A2(new_n966), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n509), .A2(new_n968), .A3(new_n513), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n970), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1971), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n509), .A2(new_n513), .A3(new_n1006), .A4(new_n968), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1008));
  AND4_X1   g583(.A1(new_n804), .A2(new_n967), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1001), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT115), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1000), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n509), .A2(new_n513), .A3(KEYINPUT45), .A4(new_n968), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n967), .A2(new_n1015), .A3(new_n971), .ZN(new_n1016));
  INV_X1    g591(.A(G1966), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n958), .A2(new_n966), .B1(new_n987), .B2(new_n1006), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n757), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1001), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G168), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1014), .A2(KEYINPUT63), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1020), .A3(new_n804), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT113), .B1(new_n1026), .B2(new_n1005), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n700), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1025), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1027), .A2(new_n1031), .A3(G8), .A4(new_n1000), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n997), .B1(new_n1024), .B2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n989), .A2(new_n991), .A3(new_n707), .ZN(new_n1035));
  INV_X1    g610(.A(new_n982), .ZN(new_n1036));
  OAI211_X1 g611(.A(G8), .B(new_n988), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1027), .A2(new_n1031), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1000), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n996), .A2(new_n1023), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT63), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(G286), .B2(G8), .ZN(new_n1047));
  NOR3_X1   g622(.A1(G168), .A2(KEYINPUT120), .A3(new_n1001), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1022), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1050), .B1(new_n1054), .B2(KEYINPUT51), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1032), .A2(new_n997), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT121), .B1(new_n1058), .B2(new_n1014), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n967), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1029), .B(new_n1011), .C1(G2090), .C2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(G8), .A3(new_n1013), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1039), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n997), .A4(new_n1032), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1028), .B2(G2078), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n785), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n972), .A2(new_n1067), .A3(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n967), .A3(new_n1015), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1057), .B1(new_n1076), .B2(KEYINPUT124), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1022), .B2(new_n1053), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1051), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1056), .B(new_n1079), .C1(new_n1080), .C2(new_n1078), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1074), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1065), .B2(new_n1059), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1043), .B1(new_n1077), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1068), .A2(G301), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT54), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n965), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1071), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1068), .A2(new_n1070), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1093), .B2(KEYINPUT122), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1068), .A2(new_n1092), .A3(new_n1095), .A4(new_n1070), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1068), .A2(new_n1092), .A3(G301), .A4(new_n1070), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT54), .B1(new_n1074), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1055), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1088), .B1(new_n1100), .B2(new_n1066), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1028), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(G299), .B(KEYINPUT57), .Z(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1060), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1348), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1069), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n967), .A2(new_n950), .A3(new_n987), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1110), .A2(new_n611), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1106), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n611), .A2(KEYINPUT119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n611), .A2(KEYINPUT119), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1125), .B(new_n1126), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT61), .B1(new_n1117), .B2(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1110), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT61), .B(new_n1109), .C1(new_n1117), .C2(KEYINPUT118), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1132));
  NAND2_X1  g707(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n988), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1103), .A2(new_n952), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1137), .B2(new_n1136), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1132), .B(new_n1134), .C1(new_n1139), .C2(new_n558), .ZN(new_n1140));
  AND4_X1   g715(.A1(KEYINPUT117), .A2(new_n1139), .A3(KEYINPUT59), .A4(new_n558), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1119), .B1(new_n1131), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1100), .A2(new_n1066), .A3(new_n1088), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1102), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n980), .B1(new_n1087), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n973), .B1(new_n951), .B2(new_n779), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT125), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n974), .A2(new_n952), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT46), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  NOR2_X1   g728(.A1(new_n727), .A2(new_n729), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n954), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n813), .A2(G2067), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n973), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1158), .A2(KEYINPUT48), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n975), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(KEYINPUT48), .B2(new_n1158), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1153), .A2(new_n1157), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT126), .B1(new_n1147), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n980), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1043), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1084), .A2(new_n1085), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1076), .A2(KEYINPUT124), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1100), .A2(new_n1066), .A3(new_n1088), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1169), .A2(new_n1101), .A3(new_n1143), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1164), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1153), .A2(new_n1157), .A3(new_n1161), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1163), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(G319), .ZN(new_n1177));
  NOR2_X1   g751(.A1(G227), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g752(.A(new_n1178), .B(KEYINPUT127), .Z(new_n1179));
  NAND4_X1  g753(.A1(new_n871), .A2(new_n660), .A3(new_n695), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n929), .A2(new_n939), .ZN(new_n1181));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1181), .ZN(G308));
  INV_X1    g756(.A(G308), .ZN(G225));
endmodule


