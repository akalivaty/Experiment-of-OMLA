

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(G2105), .A2(n523), .ZN(n879) );
  INV_X1 U552 ( .A(G2104), .ZN(n523) );
  XNOR2_X2 U553 ( .A(n529), .B(KEYINPUT66), .ZN(G160) );
  XNOR2_X1 U554 ( .A(KEYINPUT17), .B(KEYINPUT69), .ZN(n520) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  INV_X2 U556 ( .A(n745), .ZN(n761) );
  NOR2_X1 U557 ( .A1(n755), .A2(n754), .ZN(n757) );
  OR2_X1 U558 ( .A1(n745), .A2(n905), .ZN(n516) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n756) );
  BUF_X1 U560 ( .A(n613), .Z(n876) );
  XNOR2_X1 U561 ( .A(n517), .B(KEYINPUT67), .ZN(n613) );
  NOR2_X1 U562 ( .A1(n644), .A2(G651), .ZN(n649) );
  AND2_X1 U563 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U564 ( .A1(n523), .A2(G2105), .ZN(n517) );
  NAND2_X1 U565 ( .A1(G125), .A2(n613), .ZN(n518) );
  XNOR2_X1 U566 ( .A(n518), .B(KEYINPUT68), .ZN(n528) );
  XNOR2_X2 U567 ( .A(n520), .B(n519), .ZN(n880) );
  NAND2_X1 U568 ( .A1(G137), .A2(n880), .ZN(n522) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  NAND2_X1 U570 ( .A1(G113), .A2(n875), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n526) );
  NAND2_X1 U572 ( .A1(G101), .A2(n879), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT23), .B(n524), .ZN(n525) );
  NOR2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n650) );
  NAND2_X1 U576 ( .A1(G89), .A2(n650), .ZN(n530) );
  XNOR2_X1 U577 ( .A(n530), .B(KEYINPUT4), .ZN(n531) );
  XNOR2_X1 U578 ( .A(n531), .B(KEYINPUT78), .ZN(n533) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  INV_X1 U580 ( .A(G651), .ZN(n535) );
  NOR2_X1 U581 ( .A1(n644), .A2(n535), .ZN(n651) );
  NAND2_X1 U582 ( .A1(G76), .A2(n651), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n534), .B(KEYINPUT5), .ZN(n541) );
  NOR2_X1 U585 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n536), .Z(n654) );
  NAND2_X1 U587 ( .A1(G63), .A2(n654), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G51), .A2(n649), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U592 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U593 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U594 ( .A1(G102), .A2(n879), .ZN(n544) );
  NAND2_X1 U595 ( .A1(G138), .A2(n880), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G114), .A2(n875), .ZN(n546) );
  NAND2_X1 U598 ( .A1(G126), .A2(n613), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U600 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U601 ( .A1(G85), .A2(n650), .ZN(n550) );
  NAND2_X1 U602 ( .A1(G72), .A2(n651), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U604 ( .A1(G60), .A2(n654), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G47), .A2(n649), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U607 ( .A1(n554), .A2(n553), .ZN(G290) );
  XOR2_X1 U608 ( .A(G2443), .B(G2446), .Z(n556) );
  XNOR2_X1 U609 ( .A(G2427), .B(G2451), .ZN(n555) );
  XNOR2_X1 U610 ( .A(n556), .B(n555), .ZN(n562) );
  XOR2_X1 U611 ( .A(G2430), .B(G2454), .Z(n558) );
  XNOR2_X1 U612 ( .A(G1341), .B(G1348), .ZN(n557) );
  XNOR2_X1 U613 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U614 ( .A(G2435), .B(G2438), .Z(n559) );
  XNOR2_X1 U615 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U616 ( .A(n562), .B(n561), .Z(n563) );
  AND2_X1 U617 ( .A1(G14), .A2(n563), .ZN(G401) );
  NAND2_X1 U618 ( .A1(G64), .A2(n654), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G52), .A2(n649), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U621 ( .A1(G90), .A2(n650), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G77), .A2(n651), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U625 ( .A1(n570), .A2(n569), .ZN(G171) );
  AND2_X1 U626 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U627 ( .A(G108), .ZN(G238) );
  XOR2_X1 U628 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n572) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U630 ( .A(n572), .B(n571), .ZN(G223) );
  INV_X1 U631 ( .A(G567), .ZN(n685) );
  NOR2_X1 U632 ( .A1(n685), .A2(G223), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U634 ( .A1(n650), .A2(G81), .ZN(n574) );
  XNOR2_X1 U635 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G68), .A2(n651), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n577) );
  XNOR2_X1 U639 ( .A(n578), .B(n577), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n654), .A2(G56), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n579), .Z(n580) );
  NOR2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n649), .A2(G43), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n960) );
  INV_X1 U645 ( .A(G860), .ZN(n824) );
  OR2_X1 U646 ( .A1(n960), .A2(n824), .ZN(G153) );
  XNOR2_X1 U647 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(KEYINPUT76), .ZN(n594) );
  NAND2_X1 U650 ( .A1(G79), .A2(n651), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G54), .A2(n649), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G92), .A2(n650), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G66), .A2(n654), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT77), .B(n589), .Z(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n592), .Z(n978) );
  OR2_X1 U659 ( .A1(G868), .A2(n978), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U661 ( .A1(n654), .A2(G65), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n595), .B(KEYINPUT70), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G53), .A2(n649), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U665 ( .A(KEYINPUT71), .B(n598), .ZN(n602) );
  NAND2_X1 U666 ( .A1(G91), .A2(n650), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G78), .A2(n651), .ZN(n599) );
  AND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(G299) );
  INV_X1 U670 ( .A(G868), .ZN(n668) );
  NOR2_X1 U671 ( .A1(G286), .A2(n668), .ZN(n604) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n824), .A2(G559), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n605), .A2(n978), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G559), .A2(n668), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n978), .A2(n607), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT79), .ZN(n610) );
  NOR2_X1 U680 ( .A1(n960), .A2(G868), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n879), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G111), .A2(n875), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n621) );
  XOR2_X1 U685 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n615) );
  NAND2_X1 U686 ( .A1(G123), .A2(n876), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n880), .A2(G135), .ZN(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT81), .B(n616), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U691 ( .A(KEYINPUT82), .B(n619), .Z(n620) );
  NOR2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n937) );
  XNOR2_X1 U693 ( .A(n937), .B(G2096), .ZN(n623) );
  INV_X1 U694 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G75), .A2(n651), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n624), .B(KEYINPUT88), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G50), .A2(n649), .ZN(n625) );
  XOR2_X1 U699 ( .A(KEYINPUT87), .B(n625), .Z(n626) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G88), .A2(n650), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G62), .A2(n654), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(G166) );
  NAND2_X1 U705 ( .A1(G86), .A2(n650), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G61), .A2(n654), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n651), .A2(G73), .ZN(n634) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n649), .A2(G48), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G49), .A2(n649), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U716 ( .A(KEYINPUT85), .B(n641), .Z(n642) );
  NOR2_X1 U717 ( .A1(n654), .A2(n642), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(KEYINPUT86), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n644), .A2(G87), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(G288) );
  XNOR2_X1 U721 ( .A(G166), .B(G299), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n647), .B(G305), .ZN(n648) );
  XNOR2_X1 U723 ( .A(KEYINPUT19), .B(n648), .ZN(n662) );
  NAND2_X1 U724 ( .A1(G55), .A2(n649), .ZN(n659) );
  NAND2_X1 U725 ( .A1(G93), .A2(n650), .ZN(n653) );
  NAND2_X1 U726 ( .A1(G80), .A2(n651), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U728 ( .A1(G67), .A2(n654), .ZN(n655) );
  XNOR2_X1 U729 ( .A(KEYINPUT83), .B(n655), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(KEYINPUT84), .ZN(n825) );
  XNOR2_X1 U733 ( .A(G290), .B(n825), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(G288), .ZN(n891) );
  NAND2_X1 U736 ( .A1(G559), .A2(n978), .ZN(n664) );
  XOR2_X1 U737 ( .A(n960), .B(n664), .Z(n823) );
  XNOR2_X1 U738 ( .A(n891), .B(n823), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT89), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n666), .A2(G868), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n667), .B(KEYINPUT90), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n825), .A2(n668), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U750 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n676) );
  NAND2_X1 U752 ( .A1(G132), .A2(G82), .ZN(n675) );
  XNOR2_X1 U753 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U754 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G96), .A2(n678), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT92), .B(n679), .Z(n827) );
  INV_X1 U757 ( .A(n827), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n680), .A2(G2106), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT93), .ZN(n687) );
  NAND2_X1 U760 ( .A1(G69), .A2(G120), .ZN(n682) );
  NOR2_X1 U761 ( .A1(G237), .A2(n682), .ZN(n683) );
  XOR2_X1 U762 ( .A(KEYINPUT94), .B(n683), .Z(n684) );
  NOR2_X1 U763 ( .A1(G238), .A2(n684), .ZN(n828) );
  NOR2_X1 U764 ( .A1(n685), .A2(n828), .ZN(n686) );
  NOR2_X1 U765 ( .A1(n687), .A2(n686), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n689) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n822) );
  NAND2_X1 U769 ( .A1(n822), .A2(G36), .ZN(G176) );
  XNOR2_X1 U770 ( .A(KEYINPUT95), .B(G166), .ZN(G303) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n690) );
  XOR2_X1 U772 ( .A(KEYINPUT65), .B(n690), .Z(n719) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n719), .A2(n721), .ZN(n813) );
  XNOR2_X1 U775 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NAND2_X1 U776 ( .A1(G104), .A2(n879), .ZN(n692) );
  NAND2_X1 U777 ( .A1(G140), .A2(n880), .ZN(n691) );
  NAND2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U779 ( .A(KEYINPUT34), .B(n693), .ZN(n698) );
  NAND2_X1 U780 ( .A1(G116), .A2(n875), .ZN(n695) );
  NAND2_X1 U781 ( .A1(G128), .A2(n876), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U783 ( .A(KEYINPUT35), .B(n696), .Z(n697) );
  NOR2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U785 ( .A(KEYINPUT36), .B(n699), .ZN(n856) );
  NOR2_X1 U786 ( .A1(n811), .A2(n856), .ZN(n941) );
  NAND2_X1 U787 ( .A1(n813), .A2(n941), .ZN(n809) );
  NAND2_X1 U788 ( .A1(G95), .A2(n879), .ZN(n701) );
  NAND2_X1 U789 ( .A1(G131), .A2(n880), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U791 ( .A(KEYINPUT96), .B(n702), .Z(n706) );
  NAND2_X1 U792 ( .A1(G107), .A2(n875), .ZN(n704) );
  NAND2_X1 U793 ( .A1(G119), .A2(n876), .ZN(n703) );
  AND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n857) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n857), .ZN(n715) );
  NAND2_X1 U797 ( .A1(G117), .A2(n875), .ZN(n708) );
  NAND2_X1 U798 ( .A1(G129), .A2(n876), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n879), .A2(G105), .ZN(n709) );
  XOR2_X1 U801 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n880), .A2(G141), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n872) );
  NAND2_X1 U805 ( .A1(G1996), .A2(n872), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n936) );
  NAND2_X1 U807 ( .A1(n936), .A2(n813), .ZN(n716) );
  XNOR2_X1 U808 ( .A(n716), .B(KEYINPUT97), .ZN(n806) );
  INV_X1 U809 ( .A(n806), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n809), .A2(n717), .ZN(n718) );
  XNOR2_X1 U811 ( .A(n718), .B(KEYINPUT98), .ZN(n801) );
  INV_X1 U812 ( .A(n719), .ZN(n720) );
  NOR2_X4 U813 ( .A1(n721), .A2(n720), .ZN(n745) );
  NAND2_X2 U814 ( .A1(G8), .A2(n761), .ZN(n794) );
  XNOR2_X1 U815 ( .A(KEYINPUT103), .B(KEYINPUT29), .ZN(n743) );
  XOR2_X1 U816 ( .A(G1996), .B(KEYINPUT101), .Z(n1000) );
  NAND2_X1 U817 ( .A1(n745), .A2(n1000), .ZN(n722) );
  XNOR2_X1 U818 ( .A(n722), .B(KEYINPUT26), .ZN(n723) );
  INV_X1 U819 ( .A(G1341), .ZN(n905) );
  NAND2_X1 U820 ( .A1(n723), .A2(n516), .ZN(n724) );
  NOR2_X1 U821 ( .A1(n960), .A2(n724), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n978), .A2(n730), .ZN(n729) );
  AND2_X1 U823 ( .A1(n745), .A2(G2067), .ZN(n725) );
  XOR2_X1 U824 ( .A(n725), .B(KEYINPUT102), .Z(n727) );
  NAND2_X1 U825 ( .A1(n761), .A2(G1348), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U827 ( .A1(n729), .A2(n728), .ZN(n732) );
  OR2_X1 U828 ( .A1(n978), .A2(n730), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n737) );
  INV_X1 U830 ( .A(G299), .ZN(n971) );
  NAND2_X1 U831 ( .A1(n745), .A2(G2072), .ZN(n733) );
  XNOR2_X1 U832 ( .A(n733), .B(KEYINPUT27), .ZN(n735) );
  XOR2_X1 U833 ( .A(KEYINPUT100), .B(G1956), .Z(n904) );
  NOR2_X1 U834 ( .A1(n745), .A2(n904), .ZN(n734) );
  NOR2_X1 U835 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U836 ( .A1(n971), .A2(n738), .ZN(n736) );
  NAND2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n741) );
  OR2_X1 U838 ( .A1(n971), .A2(n738), .ZN(n739) );
  XNOR2_X1 U839 ( .A(n739), .B(KEYINPUT28), .ZN(n740) );
  NAND2_X1 U840 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U841 ( .A(n743), .B(n742), .ZN(n749) );
  INV_X1 U842 ( .A(G1961), .ZN(n903) );
  NAND2_X1 U843 ( .A1(n761), .A2(n903), .ZN(n747) );
  XOR2_X1 U844 ( .A(G2078), .B(KEYINPUT25), .Z(n744) );
  XNOR2_X1 U845 ( .A(KEYINPUT99), .B(n744), .ZN(n994) );
  NAND2_X1 U846 ( .A1(n745), .A2(n994), .ZN(n746) );
  NAND2_X1 U847 ( .A1(n747), .A2(n746), .ZN(n753) );
  NAND2_X1 U848 ( .A1(n753), .A2(G171), .ZN(n748) );
  NAND2_X1 U849 ( .A1(n749), .A2(n748), .ZN(n759) );
  NOR2_X1 U850 ( .A1(G1966), .A2(n794), .ZN(n771) );
  NOR2_X1 U851 ( .A1(G2084), .A2(n761), .ZN(n772) );
  NOR2_X1 U852 ( .A1(n771), .A2(n772), .ZN(n750) );
  NAND2_X1 U853 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U854 ( .A(KEYINPUT30), .B(n751), .ZN(n752) );
  NOR2_X1 U855 ( .A1(n752), .A2(G168), .ZN(n755) );
  NOR2_X1 U856 ( .A1(G171), .A2(n753), .ZN(n754) );
  XNOR2_X1 U857 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U858 ( .A1(n759), .A2(n758), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n769), .A2(G286), .ZN(n766) );
  NOR2_X1 U860 ( .A1(G1971), .A2(n794), .ZN(n760) );
  XOR2_X1 U861 ( .A(KEYINPUT105), .B(n760), .Z(n763) );
  NOR2_X1 U862 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U863 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U864 ( .A1(n764), .A2(G303), .ZN(n765) );
  NAND2_X1 U865 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U866 ( .A1(G8), .A2(n767), .ZN(n768) );
  XNOR2_X1 U867 ( .A(n768), .B(KEYINPUT32), .ZN(n776) );
  XOR2_X1 U868 ( .A(KEYINPUT104), .B(n769), .Z(n770) );
  NOR2_X1 U869 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n772), .A2(G8), .ZN(n773) );
  NAND2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n792) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n782) );
  NOR2_X1 U874 ( .A1(G1971), .A2(G303), .ZN(n777) );
  NOR2_X1 U875 ( .A1(n782), .A2(n777), .ZN(n967) );
  NAND2_X1 U876 ( .A1(n792), .A2(n967), .ZN(n778) );
  NAND2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NAND2_X1 U878 ( .A1(n778), .A2(n966), .ZN(n779) );
  NOR2_X1 U879 ( .A1(n794), .A2(n779), .ZN(n780) );
  XNOR2_X1 U880 ( .A(n780), .B(KEYINPUT64), .ZN(n781) );
  NOR2_X1 U881 ( .A1(n781), .A2(KEYINPUT33), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n782), .A2(KEYINPUT33), .ZN(n783) );
  NOR2_X1 U883 ( .A1(n783), .A2(n794), .ZN(n784) );
  NOR2_X1 U884 ( .A1(n785), .A2(n784), .ZN(n787) );
  XOR2_X1 U885 ( .A(G1981), .B(KEYINPUT106), .Z(n786) );
  XNOR2_X1 U886 ( .A(G305), .B(n786), .ZN(n963) );
  NAND2_X1 U887 ( .A1(n787), .A2(n963), .ZN(n799) );
  NOR2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XOR2_X1 U889 ( .A(n788), .B(KEYINPUT24), .Z(n789) );
  OR2_X1 U890 ( .A1(n794), .A2(n789), .ZN(n797) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n790) );
  XOR2_X1 U892 ( .A(KEYINPUT107), .B(n790), .Z(n791) );
  NAND2_X1 U893 ( .A1(G8), .A2(n791), .ZN(n793) );
  NAND2_X1 U894 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n795), .A2(n794), .ZN(n796) );
  AND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n803) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n976) );
  NAND2_X1 U900 ( .A1(n976), .A2(n813), .ZN(n802) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n816) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n872), .ZN(n932) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n857), .ZN(n935) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U905 ( .A1(n935), .A2(n804), .ZN(n805) );
  NOR2_X1 U906 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n932), .A2(n807), .ZN(n808) );
  XNOR2_X1 U908 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n811), .A2(n856), .ZN(n945) );
  NAND2_X1 U911 ( .A1(n812), .A2(n945), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U914 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n818), .B(n817), .ZN(G329) );
  INV_X1 U916 ( .A(G223), .ZN(n819) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U919 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U921 ( .A1(n822), .A2(n821), .ZN(G188) );
  NAND2_X1 U923 ( .A1(n824), .A2(n823), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n826), .B(n825), .ZN(G145) );
  INV_X1 U925 ( .A(G132), .ZN(G219) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(G82), .ZN(G220) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NAND2_X1 U930 ( .A1(n828), .A2(n827), .ZN(G261) );
  INV_X1 U931 ( .A(G261), .ZN(G325) );
  XOR2_X1 U932 ( .A(G2100), .B(G2096), .Z(n830) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(G2678), .ZN(n829) );
  XNOR2_X1 U934 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U935 ( .A(KEYINPUT43), .B(G2090), .Z(n832) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U937 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U938 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U939 ( .A(G2084), .B(G2078), .ZN(n835) );
  XNOR2_X1 U940 ( .A(n836), .B(n835), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1981), .B(G1971), .Z(n838) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1961), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U944 ( .A(G1976), .B(G1966), .Z(n840) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U946 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U947 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U948 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n843) );
  XNOR2_X1 U949 ( .A(n844), .B(n843), .ZN(n846) );
  XOR2_X1 U950 ( .A(G1956), .B(G2474), .Z(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G124), .A2(n876), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n847), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U954 ( .A1(G100), .A2(n879), .ZN(n848) );
  XOR2_X1 U955 ( .A(KEYINPUT111), .B(n848), .Z(n849) );
  NAND2_X1 U956 ( .A1(n850), .A2(n849), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n880), .A2(G136), .ZN(n851) );
  XNOR2_X1 U958 ( .A(n851), .B(KEYINPUT110), .ZN(n853) );
  NAND2_X1 U959 ( .A1(G112), .A2(n875), .ZN(n852) );
  NAND2_X1 U960 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U961 ( .A1(n855), .A2(n854), .ZN(G162) );
  XNOR2_X1 U962 ( .A(G164), .B(n856), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U964 ( .A(n859), .B(KEYINPUT114), .Z(n861) );
  XNOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U967 ( .A(G162), .B(n862), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G103), .A2(n879), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G139), .A2(n880), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n875), .A2(G115), .ZN(n865) );
  XNOR2_X1 U972 ( .A(n865), .B(KEYINPUT112), .ZN(n867) );
  NAND2_X1 U973 ( .A1(G127), .A2(n876), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U977 ( .A(KEYINPUT113), .B(n871), .Z(n947) );
  XNOR2_X1 U978 ( .A(n872), .B(n947), .ZN(n873) );
  XNOR2_X1 U979 ( .A(n874), .B(n873), .ZN(n889) );
  NAND2_X1 U980 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G142), .A2(n880), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n886), .B(G160), .ZN(n887) );
  XOR2_X1 U989 ( .A(n937), .B(n887), .Z(n888) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U991 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n960), .B(G171), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(n978), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(G37), .A2(n895), .ZN(n896) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n896), .Z(G397) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n897) );
  XOR2_X1 U999 ( .A(KEYINPUT49), .B(n897), .Z(n898) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n898), .ZN(n899) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n899), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(n900), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1006 ( .A(G5), .B(n903), .ZN(n924) );
  XNOR2_X1 U1007 ( .A(n904), .B(G20), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n905), .B(G19), .ZN(n908) );
  XOR2_X1 U1009 ( .A(G1981), .B(G6), .Z(n906) );
  XNOR2_X1 U1010 ( .A(KEYINPUT126), .B(n906), .ZN(n907) );
  NAND2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n911) );
  XOR2_X1 U1012 ( .A(KEYINPUT59), .B(G1348), .Z(n909) );
  XNOR2_X1 U1013 ( .A(G4), .B(n909), .ZN(n910) );
  NOR2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(n914), .B(KEYINPUT60), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(G1986), .B(G24), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(G22), .B(G1971), .ZN(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G1976), .B(KEYINPUT127), .ZN(n917) );
  XNOR2_X1 U1021 ( .A(n917), .B(G23), .ZN(n918) );
  NAND2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(KEYINPUT58), .B(n920), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G21), .B(G1966), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT61), .B(n927), .ZN(n929) );
  INV_X1 U1029 ( .A(G16), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n930), .A2(G11), .ZN(n959) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n933), .Z(n943) );
  XOR2_X1 U1035 ( .A(G2084), .B(G160), .Z(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(KEYINPUT117), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1043 ( .A(G2072), .B(n947), .Z(n949) );
  XOR2_X1 U1044 ( .A(G164), .B(G2078), .Z(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1046 ( .A(KEYINPUT50), .B(n950), .Z(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n953), .ZN(n955) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G29), .ZN(n957) );
  XOR2_X1 U1052 ( .A(KEYINPUT118), .B(n957), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n989) );
  XNOR2_X1 U1054 ( .A(G16), .B(KEYINPUT56), .ZN(n987) );
  XOR2_X1 U1055 ( .A(n960), .B(G1341), .Z(n962) );
  XNOR2_X1 U1056 ( .A(G171), .B(G1961), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n984) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT57), .ZN(n982) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n969) );
  AND2_X1 U1062 ( .A1(G303), .A2(G1971), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1064 ( .A(KEYINPUT122), .B(n970), .Z(n973) );
  XOR2_X1 U1065 ( .A(n971), .B(G1956), .Z(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT123), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT124), .B(n977), .Z(n980) );
  XOR2_X1 U1070 ( .A(n978), .B(G1348), .Z(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n1013) );
  XNOR2_X1 U1077 ( .A(KEYINPUT119), .B(G2067), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n990), .B(G26), .ZN(n999) );
  XNOR2_X1 U1079 ( .A(G1991), .B(G25), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G33), .B(G2072), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(G28), .A2(n993), .ZN(n997) );
  XOR2_X1 U1083 ( .A(G27), .B(n994), .Z(n995) );
  XNOR2_X1 U1084 ( .A(KEYINPUT120), .B(n995), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XOR2_X1 U1087 ( .A(G32), .B(n1000), .Z(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT121), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1090 ( .A(KEYINPUT53), .B(n1004), .Z(n1007) );
  XOR2_X1 U1091 ( .A(G34), .B(KEYINPUT54), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(G2084), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G35), .B(G2090), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(KEYINPUT55), .B(n1010), .Z(n1011) );
  NOR2_X1 U1097 ( .A1(G29), .A2(n1011), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

