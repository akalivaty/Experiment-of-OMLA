//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G15gat), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G1gat), .ZN(new_n212));
  OAI21_X1  g011(.A(G8gat), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT88), .B1(new_n211), .B2(new_n207), .ZN(new_n215));
  INV_X1    g014(.A(G8gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(new_n205), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n213), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n214), .B1(new_n213), .B2(new_n219), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G43gat), .A2(G50gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT15), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  INV_X1    g026(.A(G29gat), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G43gat), .ZN(new_n233));
  INV_X1    g032(.A(G50gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT15), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n223), .ZN(new_n237));
  NAND2_X1  g036(.A1(G29gat), .A2(G36gat), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n226), .A2(new_n232), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT86), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n230), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n243), .A2(new_n238), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n239), .B1(new_n244), .B2(new_n226), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT90), .B1(new_n222), .B2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n210), .A2(new_n212), .A3(G8gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n216), .B1(new_n215), .B2(new_n218), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT89), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n213), .A2(new_n219), .A3(new_n214), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n226), .B1(new_n243), .B2(new_n238), .ZN(new_n255));
  AND4_X1   g054(.A1(new_n226), .A2(new_n232), .A3(new_n237), .A4(new_n238), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT92), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n259));
  AOI211_X1 g058(.A(new_n259), .B(new_n245), .C1(new_n249), .C2(new_n250), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n246), .A2(new_n253), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G229gat), .A2(G233gat), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT13), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT17), .B1(new_n245), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n265), .B(KEYINPUT17), .C1(new_n255), .C2(new_n256), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n213), .B(new_n219), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n262), .B(new_n269), .C1(new_n246), .C2(new_n253), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT18), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n251), .B(new_n252), .ZN(new_n274));
  INV_X1    g073(.A(new_n272), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n274), .A2(new_n262), .A3(new_n269), .A4(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n264), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G141gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT11), .ZN(new_n279));
  INV_X1    g078(.A(G169gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G197gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT12), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n264), .A2(new_n283), .A3(new_n273), .A4(new_n276), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n298), .B2(new_n295), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n289), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT64), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n289), .C1(new_n294), .C2(new_n299), .ZN(new_n303));
  INV_X1    g102(.A(new_n299), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT65), .B(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT25), .B(new_n304), .C1(new_n307), .C2(new_n292), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n301), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT27), .B(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT28), .Z(new_n312));
  INV_X1    g111(.A(new_n295), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT66), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n280), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n319), .B2(new_n313), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n315), .B1(new_n320), .B2(new_n314), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n321), .A3(new_n290), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n309), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT72), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n324), .A2(new_n328), .B1(new_n325), .B2(new_n323), .ZN(new_n329));
  XNOR2_X1  g128(.A(G197gat), .B(G204gat), .ZN(new_n330));
  XOR2_X1   g129(.A(KEYINPUT69), .B(KEYINPUT22), .Z(new_n331));
  INV_X1    g130(.A(G211gat), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n335), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT71), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n326), .B1(new_n323), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n324), .B2(new_n325), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n323), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n326), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n343), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n341), .B1(new_n349), .B2(new_n340), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n354), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n345), .A2(new_n348), .ZN(new_n357));
  INV_X1    g156(.A(new_n343), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n339), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n360), .B2(new_n341), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT74), .B1(new_n350), .B2(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n360), .A2(new_n364), .A3(new_n341), .A4(new_n356), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n365), .A3(new_n351), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT35), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n370));
  INV_X1    g169(.A(G155gat), .ZN(new_n371));
  INV_X1    g170(.A(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  XOR2_X1   g173(.A(G141gat), .B(G148gat), .Z(new_n375));
  AOI211_X1 g174(.A(new_n373), .B(new_n374), .C1(new_n375), .C2(KEYINPUT75), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n377), .B2(new_n373), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n376), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n381));
  INV_X1    g180(.A(G127gat), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n382), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT67), .ZN(new_n385));
  XNOR2_X1  g184(.A(G113gat), .B(G120gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT68), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n387), .B2(KEYINPUT1), .ZN(new_n388));
  INV_X1    g187(.A(new_n386), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT76), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n379), .A2(new_n393), .A3(KEYINPUT3), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n376), .A2(new_n378), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n378), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n381), .A2(new_n392), .A3(new_n394), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  OR3_X1    g199(.A1(new_n379), .A2(new_n392), .A3(KEYINPUT4), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT4), .B1(new_n379), .B2(new_n392), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n379), .A2(new_n392), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT77), .ZN(new_n406));
  INV_X1    g205(.A(new_n379), .ZN(new_n407));
  INV_X1    g206(.A(new_n392), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n400), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT5), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n399), .A2(new_n403), .ZN(new_n413));
  INV_X1    g212(.A(new_n400), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT78), .ZN(new_n419));
  XOR2_X1   g218(.A(G57gat), .B(G85gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n370), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n411), .A2(new_n421), .A3(new_n415), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n411), .A2(new_n421), .A3(new_n415), .A4(new_n370), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n323), .A2(new_n408), .ZN(new_n428));
  INV_X1    g227(.A(G227gat), .ZN(new_n429));
  INV_X1    g228(.A(G233gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n309), .A2(new_n392), .A3(new_n322), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT32), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n433), .B(KEYINPUT32), .C1(new_n435), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n432), .ZN(new_n445));
  INV_X1    g244(.A(new_n431), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI211_X1 g246(.A(KEYINPUT34), .B(new_n431), .C1(new_n428), .C2(new_n432), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n440), .A3(new_n442), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n338), .A2(KEYINPUT29), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n396), .B1(new_n455), .B2(KEYINPUT81), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n379), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n398), .A2(new_n342), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n339), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n458), .A2(G228gat), .A3(G233gat), .A4(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n335), .B(new_n336), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n396), .B1(new_n462), .B2(KEYINPUT29), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n379), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G228gat), .A2(G233gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n461), .A2(new_n467), .A3(new_n202), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n202), .B1(new_n461), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n454), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G22gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n461), .A2(new_n467), .A3(new_n202), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n453), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(new_n234), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n470), .A2(new_n474), .A3(new_n477), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n452), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n368), .A2(new_n369), .A3(new_n427), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n362), .A2(new_n366), .A3(new_n427), .ZN(new_n483));
  INV_X1    g282(.A(new_n481), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT35), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n470), .A2(new_n474), .A3(new_n477), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n477), .B1(new_n470), .B2(new_n474), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT82), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n479), .A2(new_n490), .A3(new_n480), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n483), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n449), .A2(new_n495), .A3(new_n451), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n487), .A2(new_n488), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n426), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n423), .B2(new_n424), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n341), .C1(new_n349), .C2(new_n340), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n329), .B2(new_n339), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n349), .B2(new_n339), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT38), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(new_n354), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n501), .A2(new_n507), .A3(new_n363), .A4(new_n365), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n503), .A2(new_n354), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n350), .A2(KEYINPUT37), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n499), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n406), .A2(new_n400), .A3(new_n409), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n413), .A2(new_n414), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT83), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n513), .B2(new_n514), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n413), .A2(new_n520), .A3(new_n414), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n515), .A2(new_n517), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n413), .B2(new_n414), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n525), .A3(new_n422), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT40), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n528), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n522), .A2(new_n525), .A3(new_n422), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n424), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n366), .B2(new_n362), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n493), .B(new_n497), .C1(new_n512), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n288), .B1(new_n486), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(KEYINPUT96), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT9), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G57gat), .ZN(new_n543));
  INV_X1    g342(.A(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G57gat), .A2(G64gat), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT94), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n548), .B2(new_n549), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n555), .A2(new_n556), .A3(new_n550), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n555), .B2(new_n550), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT21), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n554), .B(KEYINPUT95), .C1(new_n557), .C2(new_n558), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n569));
  AND3_X1   g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n567), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n539), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n568), .ZN(new_n573));
  INV_X1    g372(.A(new_n569), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n538), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n561), .ZN(new_n578));
  INV_X1    g377(.A(new_n563), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT21), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n254), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n572), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n572), .B2(new_n577), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n536), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n581), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n570), .A2(new_n571), .A3(new_n539), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n538), .B1(new_n575), .B2(new_n576), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n577), .A3(new_n581), .ZN(new_n589));
  INV_X1    g388(.A(new_n536), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G99gat), .B(G106gat), .Z(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n606), .A2(new_n245), .B1(KEYINPUT41), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n605), .B1(new_n266), .B2(new_n268), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT98), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n257), .B2(KEYINPUT87), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n267), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n605), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n610), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n593), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n616), .B1(new_n615), .B2(new_n605), .ZN(new_n622));
  AOI211_X1 g421(.A(KEYINPUT98), .B(new_n606), .C1(new_n614), .C2(new_n267), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n609), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(KEYINPUT99), .A3(new_n619), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n620), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n621), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT97), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n634), .A3(new_n631), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n592), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n561), .A2(new_n563), .A3(new_n605), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n557), .A2(new_n558), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n601), .B2(new_n602), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n604), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n601), .A2(new_n642), .A3(new_n602), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n641), .A2(new_n644), .A3(new_n554), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n639), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI211_X1 g449(.A(KEYINPUT101), .B(new_n648), .C1(new_n640), .C2(new_n646), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n640), .A2(new_n654), .A3(new_n646), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n605), .A2(new_n654), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n578), .B2(new_n579), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n658), .B2(new_n648), .ZN(new_n659));
  AOI211_X1 g458(.A(KEYINPUT102), .B(new_n649), .C1(new_n655), .C2(new_n657), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n652), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(KEYINPUT103), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n658), .A2(new_n648), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT103), .B1(new_n661), .B2(new_n664), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n638), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n535), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n427), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n206), .ZN(G1324gat));
  AND2_X1   g475(.A1(new_n535), .A2(new_n673), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n367), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT42), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n674), .B2(new_n368), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(KEYINPUT42), .A3(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n680), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n452), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n677), .A2(new_n204), .A3(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n494), .A2(KEYINPUT105), .A3(new_n496), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n494), .B2(new_n496), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n674), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(G1326gat));
  INV_X1    g492(.A(new_n492), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n636), .A2(new_n637), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n582), .A2(new_n583), .A3(new_n536), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n590), .B1(new_n588), .B2(new_n589), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n671), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n535), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(G29gat), .A3(new_n427), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT45), .Z(new_n706));
  OAI211_X1 g505(.A(new_n493), .B(new_n691), .C1(new_n512), .C2(new_n533), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n486), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n698), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n486), .B2(new_n534), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n702), .A2(new_n701), .A3(new_n288), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT106), .B1(new_n715), .B2(new_n427), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n715), .A2(KEYINPUT106), .A3(new_n427), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n706), .B1(new_n717), .B2(new_n718), .ZN(G1328gat));
  NAND4_X1  g518(.A1(new_n535), .A2(new_n229), .A3(new_n367), .A4(new_n703), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT107), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n715), .B2(new_n368), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n721), .A2(new_n724), .A3(KEYINPUT46), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n722), .B(new_n723), .C1(new_n725), .C2(new_n726), .ZN(G1329gat));
  OAI21_X1  g526(.A(new_n233), .B1(new_n704), .B2(new_n452), .ZN(new_n728));
  INV_X1    g527(.A(new_n691), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n715), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n715), .B2(new_n499), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n704), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n694), .A2(G50gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n737), .A3(KEYINPUT48), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n713), .A2(new_n492), .A3(new_n714), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n735), .A2(new_n736), .B1(new_n739), .B2(G50gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g540(.A1(new_n630), .A2(new_n634), .A3(new_n631), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n634), .B1(new_n630), .B2(new_n631), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n701), .B(new_n288), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n671), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n708), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n427), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n543), .ZN(G1332gat));
  INV_X1    g547(.A(new_n746), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n367), .B1(new_n750), .B2(new_n544), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT110), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n544), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1333gat));
  AOI21_X1  g554(.A(G71gat), .B1(new_n749), .B2(new_n687), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n749), .A2(G71gat), .A3(new_n729), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(KEYINPUT111), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(KEYINPUT111), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n758), .B2(new_n759), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n749), .A2(new_n492), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n701), .A2(new_n287), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n671), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n698), .B1(new_n486), .B2(new_n707), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n486), .A2(new_n534), .ZN(new_n770));
  OAI221_X1 g569(.A(new_n768), .B1(new_n769), .B2(KEYINPUT44), .C1(new_n770), .C2(new_n711), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n427), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n769), .B2(new_n766), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n702), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n501), .A2(new_n595), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  NOR3_X1   g576(.A1(new_n368), .A2(G92gat), .A3(new_n671), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n773), .B2(new_n774), .ZN(new_n779));
  INV_X1    g578(.A(new_n768), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n710), .A2(new_n368), .A3(new_n712), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n596), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n781), .B2(new_n596), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI221_X1 g585(.A(new_n779), .B1(new_n783), .B2(KEYINPUT52), .C1(new_n781), .C2(new_n596), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n771), .B2(new_n691), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n452), .A2(G99gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n775), .B2(new_n790), .ZN(G1338gat));
  OAI21_X1  g590(.A(G106gat), .B1(new_n771), .B2(new_n499), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n499), .A2(G106gat), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n702), .B(new_n794), .C1(new_n773), .C2(new_n774), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G106gat), .B1(new_n771), .B2(new_n694), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n793), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n261), .A2(new_n263), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n262), .B1(new_n274), .B2(new_n269), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n282), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n286), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n669), .B2(new_n670), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT54), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n655), .A2(new_n649), .A3(new_n657), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n667), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n664), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n658), .A2(new_n653), .A3(new_n648), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n664), .A4(new_n809), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n287), .A2(new_n811), .A3(new_n668), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n805), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n817), .A3(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n698), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n811), .A2(new_n668), .A3(new_n816), .ZN(new_n823));
  OR4_X1    g622(.A1(new_n742), .A2(new_n743), .A3(new_n823), .A4(new_n803), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n592), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n744), .B2(new_n702), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n638), .A2(new_n828), .A3(new_n288), .A4(new_n671), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n694), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT116), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n367), .A2(new_n427), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n687), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n831), .B2(new_n694), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n687), .B(new_n835), .C1(new_n837), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n836), .A2(new_n841), .A3(G113gat), .A4(new_n287), .ZN(new_n842));
  INV_X1    g641(.A(G113gat), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n825), .A2(new_n592), .B1(new_n827), .B2(new_n829), .ZN(new_n844));
  INV_X1    g643(.A(new_n835), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n481), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n843), .B1(new_n847), .B2(new_n288), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n842), .A2(new_n848), .ZN(G1340gat));
  NAND4_X1  g648(.A1(new_n836), .A2(new_n841), .A3(G120gat), .A4(new_n702), .ZN(new_n850));
  INV_X1    g649(.A(G120gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n847), .B2(new_n671), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(G1341gat));
  AND3_X1   g652(.A1(new_n836), .A2(new_n841), .A3(new_n701), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n701), .A2(new_n382), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n854), .A2(new_n382), .B1(new_n847), .B2(new_n855), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n836), .A2(new_n841), .A3(new_n709), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G134gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n368), .A2(new_n709), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT118), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n844), .A2(new_n427), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n484), .A2(G134gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT56), .Z(new_n865));
  NAND2_X1  g664(.A1(new_n858), .A2(new_n865), .ZN(G1343gat));
  NOR2_X1   g665(.A1(new_n729), .A2(new_n499), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n846), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(G141gat), .A3(new_n288), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n694), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n805), .A2(KEYINPUT119), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n804), .B(new_n873), .C1(new_n669), .C2(new_n670), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n823), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n811), .A2(new_n816), .A3(KEYINPUT120), .A4(new_n668), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n288), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n698), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n701), .B1(new_n880), .B2(new_n824), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n827), .A2(new_n829), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT121), .B(new_n871), .C1(new_n881), .C2(new_n882), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n870), .B1(new_n844), .B2(new_n499), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n845), .A2(new_n729), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n287), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n869), .B1(new_n890), .B2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(new_n869), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n897), .B2(KEYINPUT58), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n891), .A2(KEYINPUT122), .A3(new_n892), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(G1344gat));
  AND2_X1   g699(.A1(new_n862), .A2(new_n867), .ZN(new_n901));
  INV_X1    g700(.A(G148gat), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n368), .A4(new_n702), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT123), .Z(new_n904));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n902), .C1(new_n905), .C2(new_n702), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n870), .B1(new_n831), .B2(new_n498), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n744), .A2(new_n702), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n881), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n492), .A2(new_n870), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n702), .A3(new_n889), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n904), .B1(new_n906), .B2(new_n915), .ZN(G1345gat));
  NOR2_X1   g715(.A1(new_n868), .A2(new_n592), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  AOI21_X1  g717(.A(G155gat), .B1(new_n917), .B2(KEYINPUT124), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n592), .A2(new_n371), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n918), .A2(new_n919), .B1(new_n905), .B2(new_n920), .ZN(G1346gat));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n372), .A3(new_n861), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n905), .A2(new_n709), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n372), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n368), .A2(new_n501), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n687), .B(new_n925), .C1(new_n837), .C2(new_n839), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n280), .A3(new_n288), .ZN(new_n927));
  INV_X1    g726(.A(new_n925), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n844), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n481), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n287), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n927), .A2(new_n932), .ZN(G1348gat));
  OAI21_X1  g732(.A(G176gat), .B1(new_n926), .B2(new_n671), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n318), .A3(new_n702), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  OAI21_X1  g735(.A(G183gat), .B1(new_n926), .B2(new_n592), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n310), .A3(new_n701), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT60), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n931), .A2(new_n305), .A3(new_n709), .ZN(new_n944));
  OAI21_X1  g743(.A(G190gat), .B1(new_n926), .B2(new_n698), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT61), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n947), .B(G190gat), .C1(new_n926), .C2(new_n698), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(new_n946), .B2(new_n949), .ZN(G1351gat));
  AND2_X1   g749(.A1(new_n929), .A2(new_n867), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n287), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n928), .A2(new_n729), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n844), .A2(new_n499), .ZN(new_n954));
  OAI221_X1 g753(.A(new_n953), .B1(new_n910), .B2(new_n911), .C1(new_n954), .C2(new_n870), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n287), .A2(G197gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  NOR2_X1   g757(.A1(new_n671), .A2(G204gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n929), .A2(new_n867), .A3(new_n959), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT62), .Z(new_n961));
  NAND3_X1  g760(.A1(new_n913), .A2(new_n702), .A3(new_n953), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G204gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT125), .ZN(G1353gat));
  NAND3_X1  g764(.A1(new_n951), .A2(new_n332), .A3(new_n701), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n913), .A2(new_n967), .A3(new_n701), .A4(new_n953), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(new_n955), .B2(new_n592), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND4_X1   g770(.A1(KEYINPUT63), .A2(new_n970), .A3(new_n968), .A4(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n955), .B2(new_n698), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n951), .A2(new_n333), .A3(new_n709), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n976), .B(KEYINPUT127), .Z(G1355gat));
endmodule


