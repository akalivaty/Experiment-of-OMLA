

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n825), .A2(n768), .ZN(n521) );
  BUF_X1 U554 ( .A(n704), .Z(n726) );
  OR2_X1 U555 ( .A1(n710), .A2(n709), .ZN(n722) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n723) );
  NOR2_X1 U557 ( .A1(n694), .A2(n785), .ZN(n704) );
  INV_X1 U558 ( .A(n704), .ZN(n742) );
  NOR2_X1 U559 ( .A1(G164), .A2(G1384), .ZN(n786) );
  NOR2_X1 U560 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U561 ( .A1(G651), .A2(n651), .ZN(n661) );
  AND2_X1 U562 ( .A1(n541), .A2(G2104), .ZN(n883) );
  NOR2_X2 U563 ( .A1(G2104), .A2(n541), .ZN(n886) );
  NOR2_X1 U564 ( .A1(n547), .A2(n546), .ZN(G160) );
  INV_X1 U565 ( .A(G651), .ZN(n530) );
  NOR2_X1 U566 ( .A1(G543), .A2(n530), .ZN(n522) );
  XOR2_X1 U567 ( .A(KEYINPUT1), .B(n522), .Z(n664) );
  NAND2_X1 U568 ( .A1(n664), .A2(G63), .ZN(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(KEYINPUT78), .ZN(n526) );
  XNOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT66), .B(n524), .Z(n651) );
  NAND2_X1 U572 ( .A1(G51), .A2(n661), .ZN(n525) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U574 ( .A(KEYINPUT6), .B(n527), .ZN(n535) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n660) );
  NAND2_X1 U576 ( .A1(G89), .A2(n660), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT4), .B(n528), .Z(n529) );
  XNOR2_X1 U578 ( .A(n529), .B(KEYINPUT77), .ZN(n532) );
  NOR2_X2 U579 ( .A1(n530), .A2(n651), .ZN(n658) );
  NAND2_X1 U580 ( .A1(G76), .A2(n658), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT5), .B(n533), .Z(n534) );
  NOR2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U584 ( .A(KEYINPUT7), .B(KEYINPUT79), .ZN(n536) );
  XNOR2_X1 U585 ( .A(n537), .B(n536), .ZN(G168) );
  XOR2_X1 U586 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U588 ( .A1(n887), .A2(G113), .ZN(n540) );
  INV_X1 U589 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G101), .A2(n883), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT23), .B(n538), .Z(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n547) );
  NAND2_X1 U593 ( .A1(G125), .A2(n886), .ZN(n545) );
  XNOR2_X1 U594 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n543) );
  NOR2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n543), .B(n542), .ZN(n882) );
  NAND2_X1 U597 ( .A1(G137), .A2(n882), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n882), .A2(G138), .ZN(n550) );
  NAND2_X1 U600 ( .A1(G126), .A2(n886), .ZN(n548) );
  XOR2_X1 U601 ( .A(KEYINPUT91), .B(n548), .Z(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U603 ( .A1(G102), .A2(n883), .ZN(n552) );
  NAND2_X1 U604 ( .A1(G114), .A2(n887), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U606 ( .A1(n554), .A2(n553), .ZN(G164) );
  NAND2_X1 U607 ( .A1(n664), .A2(G64), .ZN(n555) );
  XNOR2_X1 U608 ( .A(KEYINPUT67), .B(n555), .ZN(n558) );
  NAND2_X1 U609 ( .A1(n661), .A2(G52), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT68), .B(n556), .Z(n557) );
  NOR2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U612 ( .A(KEYINPUT69), .B(n559), .ZN(n564) );
  NAND2_X1 U613 ( .A1(G90), .A2(n660), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G77), .A2(n658), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U617 ( .A1(n564), .A2(n563), .ZN(G171) );
  XOR2_X1 U618 ( .A(KEYINPUT108), .B(G2446), .Z(n566) );
  XNOR2_X1 U619 ( .A(G2430), .B(G2451), .ZN(n565) );
  XNOR2_X1 U620 ( .A(n566), .B(n565), .ZN(n570) );
  XOR2_X1 U621 ( .A(G2435), .B(KEYINPUT107), .Z(n568) );
  XNOR2_X1 U622 ( .A(G2438), .B(G2454), .ZN(n567) );
  XNOR2_X1 U623 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U624 ( .A(n570), .B(n569), .Z(n572) );
  XNOR2_X1 U625 ( .A(G2443), .B(G2427), .ZN(n571) );
  XNOR2_X1 U626 ( .A(n572), .B(n571), .ZN(n575) );
  XNOR2_X1 U627 ( .A(G1341), .B(KEYINPUT106), .ZN(n573) );
  XOR2_X1 U628 ( .A(n573), .B(G1348), .Z(n574) );
  XOR2_X1 U629 ( .A(n575), .B(n574), .Z(n576) );
  AND2_X1 U630 ( .A1(G14), .A2(n576), .ZN(G401) );
  INV_X1 U631 ( .A(G132), .ZN(G219) );
  INV_X1 U632 ( .A(G82), .ZN(G220) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  NAND2_X1 U634 ( .A1(G94), .A2(G452), .ZN(n577) );
  XOR2_X1 U635 ( .A(KEYINPUT70), .B(n577), .Z(G173) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U637 ( .A(n578), .B(KEYINPUT72), .ZN(n579) );
  XNOR2_X1 U638 ( .A(KEYINPUT10), .B(n579), .ZN(G223) );
  XNOR2_X1 U639 ( .A(KEYINPUT73), .B(G223), .ZN(n835) );
  NAND2_X1 U640 ( .A1(n835), .A2(G567), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U642 ( .A1(G56), .A2(n664), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n581), .Z(n587) );
  NAND2_X1 U644 ( .A1(n660), .A2(G81), .ZN(n582) );
  XNOR2_X1 U645 ( .A(n582), .B(KEYINPUT12), .ZN(n584) );
  NAND2_X1 U646 ( .A1(G68), .A2(n658), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n585), .Z(n586) );
  NOR2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n661), .A2(G43), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n978) );
  INV_X1 U652 ( .A(G860), .ZN(n614) );
  NOR2_X1 U653 ( .A1(n978), .A2(n614), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT74), .B(n590), .Z(G153) );
  INV_X1 U655 ( .A(G171), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U657 ( .A1(n658), .A2(G79), .ZN(n592) );
  INV_X1 U658 ( .A(KEYINPUT75), .ZN(n591) );
  XNOR2_X1 U659 ( .A(n592), .B(n591), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n661), .A2(G54), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n595), .B(KEYINPUT76), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G92), .A2(n660), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G66), .A2(n664), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X2 U666 ( .A(n600), .B(KEYINPUT15), .Z(n988) );
  INV_X1 U667 ( .A(n988), .ZN(n712) );
  INV_X1 U668 ( .A(G868), .ZN(n611) );
  NAND2_X1 U669 ( .A1(n712), .A2(n611), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U671 ( .A1(G91), .A2(n660), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G53), .A2(n661), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G78), .A2(n658), .ZN(n605) );
  XNOR2_X1 U675 ( .A(KEYINPUT71), .B(n605), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n664), .A2(G65), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n609), .A2(n608), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n610), .B(KEYINPUT80), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n611), .A2(G286), .ZN(n612) );
  NOR2_X1 U682 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n615), .A2(n988), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n978), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n988), .A2(G868), .ZN(n617) );
  NOR2_X1 U688 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G123), .A2(n886), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT18), .ZN(n623) );
  NAND2_X1 U692 ( .A1(G99), .A2(n883), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(n621), .Z(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G135), .A2(n882), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G111), .A2(n887), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n930) );
  XNOR2_X1 U699 ( .A(n930), .B(G2096), .ZN(n628) );
  INV_X1 U700 ( .A(G2100), .ZN(n857) );
  NAND2_X1 U701 ( .A1(n628), .A2(n857), .ZN(G156) );
  AND2_X1 U702 ( .A1(n661), .A2(G47), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G85), .A2(n660), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G72), .A2(n658), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n664), .A2(G60), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U709 ( .A1(G75), .A2(n658), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n635), .B(KEYINPUT88), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n660), .A2(G88), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G50), .A2(n661), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G62), .A2(n664), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(G166) );
  NAND2_X1 U717 ( .A1(G73), .A2(n658), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U719 ( .A1(G61), .A2(n664), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT86), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n660), .A2(G86), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G48), .A2(n661), .ZN(n646) );
  XNOR2_X1 U724 ( .A(KEYINPUT87), .B(n646), .ZN(n647) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G87), .A2(n651), .ZN(n656) );
  NAND2_X1 U728 ( .A1(G49), .A2(n661), .ZN(n653) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U731 ( .A1(n664), .A2(n654), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U733 ( .A(KEYINPUT85), .B(n657), .Z(G288) );
  NAND2_X1 U734 ( .A1(G80), .A2(n658), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(KEYINPUT82), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G93), .A2(n660), .ZN(n663) );
  NAND2_X1 U737 ( .A1(G55), .A2(n661), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U739 ( .A1(G67), .A2(n664), .ZN(n665) );
  XNOR2_X1 U740 ( .A(KEYINPUT83), .B(n665), .ZN(n666) );
  NOR2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT84), .B(n670), .Z(n841) );
  NOR2_X1 U744 ( .A1(G868), .A2(n841), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n671), .B(KEYINPUT89), .ZN(n680) );
  XNOR2_X1 U746 ( .A(KEYINPUT19), .B(G290), .ZN(n676) );
  XOR2_X1 U747 ( .A(G299), .B(G305), .Z(n672) );
  XNOR2_X1 U748 ( .A(n672), .B(n841), .ZN(n673) );
  XNOR2_X1 U749 ( .A(G166), .B(n673), .ZN(n674) );
  XNOR2_X1 U750 ( .A(n674), .B(G288), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n676), .B(n675), .ZN(n910) );
  NAND2_X1 U752 ( .A1(G559), .A2(n988), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n677), .B(n978), .ZN(n840) );
  XNOR2_X1 U754 ( .A(n910), .B(n840), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G868), .A2(n678), .ZN(n679) );
  NAND2_X1 U756 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U761 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U763 ( .A1(G120), .A2(G108), .ZN(n685) );
  NOR2_X1 U764 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G69), .A2(n686), .ZN(n844) );
  NAND2_X1 U766 ( .A1(n844), .A2(G567), .ZN(n692) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U769 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G96), .A2(n689), .ZN(n843) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n843), .ZN(n690) );
  XNOR2_X1 U772 ( .A(KEYINPUT90), .B(n690), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n692), .A2(n691), .ZN(n845) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n693) );
  NOR2_X1 U775 ( .A1(n845), .A2(n693), .ZN(n839) );
  NAND2_X1 U776 ( .A1(n839), .A2(G36), .ZN(G176) );
  XOR2_X1 U777 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  INV_X1 U778 ( .A(n786), .ZN(n694) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n785) );
  NAND2_X1 U780 ( .A1(G1996), .A2(n726), .ZN(n695) );
  XNOR2_X1 U781 ( .A(KEYINPUT26), .B(n695), .ZN(n699) );
  NAND2_X1 U782 ( .A1(G1341), .A2(n742), .ZN(n696) );
  XNOR2_X1 U783 ( .A(KEYINPUT99), .B(n696), .ZN(n697) );
  NOR2_X1 U784 ( .A1(n978), .A2(n697), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n713) );
  NOR2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(KEYINPUT100), .ZN(n710) );
  INV_X1 U788 ( .A(G1348), .ZN(n996) );
  NOR2_X1 U789 ( .A1(n726), .A2(n996), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT101), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n726), .A2(G2067), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n708) );
  INV_X1 U793 ( .A(G299), .ZN(n717) );
  NAND2_X1 U794 ( .A1(n704), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U795 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U796 ( .A(G1956), .ZN(n846) );
  NOR2_X1 U797 ( .A1(n846), .A2(n726), .ZN(n706) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n716) );
  NAND2_X1 U799 ( .A1(n717), .A2(n716), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n708), .A2(n711), .ZN(n709) );
  INV_X1 U801 ( .A(n711), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n720) );
  NOR2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U805 ( .A(n718), .B(KEYINPUT28), .Z(n719) );
  AND2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U808 ( .A(n724), .B(n723), .ZN(n731) );
  NOR2_X1 U809 ( .A1(n726), .A2(G1961), .ZN(n725) );
  XNOR2_X1 U810 ( .A(n725), .B(KEYINPUT97), .ZN(n728) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U812 ( .A1(n726), .A2(n955), .ZN(n727) );
  NAND2_X1 U813 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U814 ( .A(KEYINPUT98), .B(n729), .ZN(n735) );
  NAND2_X1 U815 ( .A1(G171), .A2(n735), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n740) );
  NAND2_X1 U817 ( .A1(G8), .A2(n742), .ZN(n825) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n825), .ZN(n755) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n742), .ZN(n752) );
  NOR2_X1 U820 ( .A1(n755), .A2(n752), .ZN(n732) );
  NAND2_X1 U821 ( .A1(G8), .A2(n732), .ZN(n733) );
  XNOR2_X1 U822 ( .A(KEYINPUT30), .B(n733), .ZN(n734) );
  NOR2_X1 U823 ( .A1(G168), .A2(n734), .ZN(n737) );
  NOR2_X1 U824 ( .A1(G171), .A2(n735), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(n738), .Z(n739) );
  NAND2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n753) );
  NAND2_X1 U828 ( .A1(n753), .A2(G286), .ZN(n741) );
  XNOR2_X1 U829 ( .A(n741), .B(KEYINPUT102), .ZN(n749) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n742), .ZN(n743) );
  XOR2_X1 U831 ( .A(KEYINPUT103), .B(n743), .Z(n745) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n825), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G303), .A2(n746), .ZN(n747) );
  XNOR2_X1 U835 ( .A(KEYINPUT104), .B(n747), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n750), .A2(G8), .ZN(n751) );
  XNOR2_X1 U838 ( .A(n751), .B(KEYINPUT32), .ZN(n817) );
  NAND2_X1 U839 ( .A1(G8), .A2(n752), .ZN(n757) );
  INV_X1 U840 ( .A(n753), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n818) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n973) );
  AND2_X1 U844 ( .A1(n818), .A2(n973), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n817), .A2(n758), .ZN(n763) );
  INV_X1 U846 ( .A(n973), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n767) );
  NOR2_X1 U848 ( .A1(G303), .A2(G1971), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n767), .A2(n759), .ZN(n982) );
  OR2_X1 U850 ( .A1(n760), .A2(n982), .ZN(n761) );
  OR2_X1 U851 ( .A1(n825), .A2(n761), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n764), .B(KEYINPUT64), .ZN(n765) );
  NOR2_X1 U854 ( .A1(KEYINPUT33), .A2(n765), .ZN(n766) );
  XNOR2_X1 U855 ( .A(n766), .B(KEYINPUT105), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n767), .A2(KEYINPUT33), .ZN(n768) );
  AND2_X1 U857 ( .A1(n769), .A2(n521), .ZN(n816) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U859 ( .A1(G105), .A2(n883), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT38), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G129), .A2(n886), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G141), .A2(n882), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n887), .A2(G117), .ZN(n773) );
  XOR2_X1 U865 ( .A(KEYINPUT96), .B(n773), .Z(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n894) );
  NOR2_X1 U868 ( .A1(G1996), .A2(n894), .ZN(n922) );
  AND2_X1 U869 ( .A1(n894), .A2(G1996), .ZN(n931) );
  NAND2_X1 U870 ( .A1(G131), .A2(n882), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G95), .A2(n883), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U873 ( .A(KEYINPUT95), .B(n780), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G119), .A2(n886), .ZN(n782) );
  NAND2_X1 U875 ( .A1(G107), .A2(n887), .ZN(n781) );
  AND2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n899) );
  AND2_X1 U878 ( .A1(n899), .A2(G1991), .ZN(n937) );
  OR2_X1 U879 ( .A1(n931), .A2(n937), .ZN(n787) );
  NOR2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n808) );
  NAND2_X1 U881 ( .A1(n787), .A2(n808), .ZN(n809) );
  INV_X1 U882 ( .A(n809), .ZN(n790) );
  NOR2_X1 U883 ( .A1(G1991), .A2(n899), .ZN(n933) );
  NOR2_X1 U884 ( .A1(G1986), .A2(G290), .ZN(n788) );
  NOR2_X1 U885 ( .A1(n933), .A2(n788), .ZN(n789) );
  NOR2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U887 ( .A1(n922), .A2(n791), .ZN(n792) );
  XNOR2_X1 U888 ( .A(n792), .B(KEYINPUT39), .ZN(n804) );
  XNOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n882), .A2(G140), .ZN(n793) );
  XOR2_X1 U891 ( .A(KEYINPUT93), .B(n793), .Z(n795) );
  NAND2_X1 U892 ( .A1(n883), .A2(G104), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(n796), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n887), .A2(G116), .ZN(n797) );
  XNOR2_X1 U896 ( .A(n797), .B(KEYINPUT94), .ZN(n799) );
  NAND2_X1 U897 ( .A1(G128), .A2(n886), .ZN(n798) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U899 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U901 ( .A(KEYINPUT36), .B(n803), .ZN(n900) );
  NOR2_X1 U902 ( .A1(n805), .A2(n900), .ZN(n941) );
  NAND2_X1 U903 ( .A1(n808), .A2(n941), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n804), .A2(n810), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n805), .A2(n900), .ZN(n942) );
  NAND2_X1 U906 ( .A1(n806), .A2(n942), .ZN(n807) );
  AND2_X1 U907 ( .A1(n807), .A2(n808), .ZN(n828) );
  INV_X1 U908 ( .A(n828), .ZN(n814) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n975) );
  AND2_X1 U910 ( .A1(n975), .A2(n808), .ZN(n812) );
  NAND2_X1 U911 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U912 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n831) );
  AND2_X1 U914 ( .A1(n983), .A2(n831), .ZN(n815) );
  NAND2_X1 U915 ( .A1(n816), .A2(n815), .ZN(n833) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n821) );
  NOR2_X1 U917 ( .A1(G2090), .A2(G303), .ZN(n819) );
  NAND2_X1 U918 ( .A1(G8), .A2(n819), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n822), .A2(n825), .ZN(n827) );
  NOR2_X1 U921 ( .A1(G1981), .A2(G305), .ZN(n823) );
  XOR2_X1 U922 ( .A(n823), .B(KEYINPUT24), .Z(n824) );
  OR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n829) );
  OR2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U928 ( .A(KEYINPUT40), .B(n834), .ZN(G329) );
  NAND2_X1 U929 ( .A1(n835), .A2(G2106), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT109), .B(n836), .Z(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  NOR2_X1 U937 ( .A1(n840), .A2(G860), .ZN(n842) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G145) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n845), .ZN(G319) );
  XOR2_X1 U944 ( .A(n846), .B(KEYINPUT41), .Z(n856) );
  XOR2_X1 U945 ( .A(G1981), .B(G1961), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U952 ( .A(KEYINPUT110), .B(G2474), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(G229) );
  XNOR2_X1 U955 ( .A(n857), .B(G2096), .ZN(n859) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(G2678), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2090), .Z(n861) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U961 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U964 ( .A1(G124), .A2(n886), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G100), .A2(n883), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT111), .B(n867), .Z(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G136), .A2(n882), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G112), .A2(n887), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G130), .A2(n886), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G118), .A2(n887), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U976 ( .A1(n883), .A2(G106), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT112), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G142), .A2(n882), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n898) );
  NAND2_X1 U982 ( .A1(G139), .A2(n882), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G103), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U985 ( .A1(G127), .A2(n886), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G115), .A2(n887), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  XNOR2_X1 U989 ( .A(KEYINPUT114), .B(n891), .ZN(n892) );
  NOR2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n924) );
  XOR2_X1 U991 ( .A(n930), .B(n924), .Z(n896) );
  XOR2_X1 U992 ( .A(G160), .B(n894), .Z(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U995 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n907) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n904) );
  XNOR2_X1 U998 ( .A(G162), .B(KEYINPUT48), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(G164), .B(n905), .Z(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1003 ( .A(G286), .B(G171), .Z(n909) );
  XNOR2_X1 U1004 ( .A(n909), .B(n978), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(n988), .B(n910), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n914) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n916), .ZN(n917) );
  XOR2_X1 U1012 ( .A(KEYINPUT115), .B(n917), .Z(n920) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(KEYINPUT116), .B(n918), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  INV_X1 U1018 ( .A(KEYINPUT55), .ZN(n946) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT51), .B(n923), .ZN(n929) );
  XOR2_X1 U1022 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT50), .B(n927), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n939) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n935) );
  XOR2_X1 U1028 ( .A(G160), .B(G2084), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1035 ( .A(KEYINPUT52), .B(n944), .Z(n945) );
  NAND2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1037 ( .A1(n947), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1038 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(n948), .B(KEYINPUT54), .ZN(n963) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1041 ( .A1(n949), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(KEYINPUT119), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G2072), .B(G33), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1047 ( .A(G2067), .B(G26), .Z(n958) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(n955), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G27), .B(n956), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(n961), .B(KEYINPUT53), .ZN(n962) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1054 ( .A(G2090), .B(KEYINPUT118), .Z(n964) );
  XNOR2_X1 U1055 ( .A(G35), .B(n964), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1057 ( .A(KEYINPUT55), .B(n967), .Z(n969) );
  INV_X1 U1058 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n970), .ZN(n1025) );
  INV_X1 U1061 ( .A(G16), .ZN(n1021) );
  XOR2_X1 U1062 ( .A(n1021), .B(KEYINPUT56), .Z(n994) );
  XOR2_X1 U1063 ( .A(G299), .B(KEYINPUT121), .Z(n971) );
  XOR2_X1 U1064 ( .A(n971), .B(G1956), .Z(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(G303), .A2(G1971), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1074 ( .A(KEYINPUT57), .B(n985), .Z(n986) );
  NOR2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n992) );
  XOR2_X1 U1076 ( .A(G171), .B(G1961), .Z(n990) );
  XOR2_X1 U1077 ( .A(n988), .B(G1348), .Z(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n1023) );
  XOR2_X1 U1081 ( .A(G1961), .B(G5), .Z(n1010) );
  XOR2_X1 U1082 ( .A(G1966), .B(G21), .Z(n995) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n995), .ZN(n1007) );
  XOR2_X1 U1084 ( .A(KEYINPUT122), .B(G4), .Z(n998) );
  XOR2_X1 U1085 ( .A(n996), .B(KEYINPUT59), .Z(n997) );
  XNOR2_X1 U1086 ( .A(n998), .B(n997), .ZN(n1004) );
  XOR2_X1 U1087 ( .A(G20), .B(G1956), .Z(n1002) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1005), .Z(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1018) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1014) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XOR2_X1 U1110 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1028) );
  XNOR2_X1 U1111 ( .A(n1029), .B(n1028), .ZN(G311) );
  XNOR2_X1 U1112 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

