

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(KEYINPUT112), .B(n531), .ZN(n542) );
  NOR2_X1 U324 ( .A1(n513), .A2(n430), .ZN(n568) );
  XNOR2_X1 U325 ( .A(n301), .B(n300), .ZN(n307) );
  NOR2_X1 U326 ( .A1(n542), .A2(n557), .ZN(n532) );
  XOR2_X1 U327 ( .A(n295), .B(n294), .Z(n291) );
  XNOR2_X1 U328 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U329 ( .A(n435), .B(n364), .ZN(n365) );
  XNOR2_X1 U330 ( .A(n296), .B(n291), .ZN(n301) );
  XNOR2_X1 U331 ( .A(n370), .B(n369), .ZN(n371) );
  INV_X1 U332 ( .A(KEYINPUT110), .ZN(n525) );
  XNOR2_X1 U333 ( .A(n372), .B(n371), .ZN(n374) );
  XNOR2_X1 U334 ( .A(n526), .B(n525), .ZN(n545) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n447) );
  XNOR2_X1 U336 ( .A(n309), .B(n308), .ZN(n554) );
  XOR2_X1 U337 ( .A(n459), .B(KEYINPUT28), .Z(n518) );
  XNOR2_X1 U338 ( .A(n447), .B(KEYINPUT58), .ZN(n448) );
  XNOR2_X1 U339 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT71), .B(KEYINPUT11), .Z(n293) );
  XNOR2_X1 U341 ( .A(G106GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n309) );
  XOR2_X1 U343 ( .A(G92GAT), .B(G85GAT), .Z(n363) );
  XNOR2_X1 U344 ( .A(G218GAT), .B(n363), .ZN(n296) );
  XOR2_X1 U345 ( .A(KEYINPUT9), .B(G134GAT), .Z(n295) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U347 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n298) );
  XNOR2_X1 U348 ( .A(G190GAT), .B(KEYINPUT65), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(n299), .B(KEYINPUT72), .Z(n300) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n302), .B(G29GAT), .ZN(n303) );
  XOR2_X1 U353 ( .A(n303), .B(KEYINPUT7), .Z(n305) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G50GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n349) );
  XNOR2_X1 U356 ( .A(n349), .B(G162GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n310), .B(KEYINPUT0), .ZN(n336) );
  XOR2_X1 U360 ( .A(n336), .B(G176GAT), .Z(n312) );
  XOR2_X1 U361 ( .A(G113GAT), .B(G169GAT), .Z(n348) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(n348), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n317) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G71GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n313), .B(G120GAT), .ZN(n366) );
  XOR2_X1 U366 ( .A(n366), .B(KEYINPUT78), .Z(n315) );
  NAND2_X1 U367 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(n317), .B(n316), .Z(n327) );
  XOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT18), .Z(n319) );
  XNOR2_X1 U371 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U373 ( .A(n320), .B(KEYINPUT80), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT17), .B(G190GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n417) );
  XOR2_X1 U376 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n324) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(KEYINPUT79), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n417), .B(n325), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n527) );
  XOR2_X1 U381 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n445) );
  XOR2_X1 U382 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n329) );
  XNOR2_X1 U383 ( .A(KEYINPUT88), .B(KEYINPUT1), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n343) );
  XOR2_X1 U385 ( .A(G57GAT), .B(G120GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G113GAT), .B(G148GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U388 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n333) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U391 ( .A(n335), .B(n334), .Z(n341) );
  XOR2_X1 U392 ( .A(G85GAT), .B(n336), .Z(n338) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(G29GAT), .B(n339), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U398 ( .A(G162GAT), .B(KEYINPUT2), .Z(n345) );
  XNOR2_X1 U399 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U401 ( .A(G155GAT), .B(n346), .Z(n431) );
  XOR2_X1 U402 ( .A(n347), .B(n431), .Z(n453) );
  INV_X1 U403 ( .A(n453), .ZN(n513) );
  XOR2_X1 U404 ( .A(KEYINPUT29), .B(n348), .Z(n351) );
  XNOR2_X1 U405 ( .A(n349), .B(G197GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U407 ( .A(KEYINPUT30), .B(G141GAT), .Z(n353) );
  NAND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n355), .B(n354), .Z(n359) );
  XOR2_X1 U411 ( .A(G1GAT), .B(G15GAT), .Z(n357) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(G22GAT), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n395) );
  XNOR2_X1 U414 ( .A(n395), .B(KEYINPUT66), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n569) );
  XOR2_X1 U416 ( .A(G78GAT), .B(G148GAT), .Z(n361) );
  XNOR2_X1 U417 ( .A(G106GAT), .B(G204GAT), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n435) );
  AND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n365), .B(KEYINPUT69), .ZN(n372) );
  XOR2_X1 U421 ( .A(n366), .B(KEYINPUT68), .Z(n370) );
  XOR2_X1 U422 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n368) );
  XNOR2_X1 U423 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n367) );
  XOR2_X1 U424 ( .A(n368), .B(n367), .Z(n369) );
  XOR2_X1 U425 ( .A(G176GAT), .B(G64GAT), .Z(n418) );
  XOR2_X1 U426 ( .A(KEYINPUT13), .B(G57GAT), .Z(n391) );
  XNOR2_X1 U427 ( .A(n418), .B(n391), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n575) );
  XNOR2_X1 U429 ( .A(n575), .B(KEYINPUT41), .ZN(n375) );
  INV_X1 U430 ( .A(n375), .ZN(n498) );
  NOR2_X1 U431 ( .A1(n569), .A2(n498), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n376), .B(KEYINPUT46), .ZN(n379) );
  INV_X1 U433 ( .A(n379), .ZN(n377) );
  NAND2_X1 U434 ( .A1(n377), .A2(KEYINPUT108), .ZN(n381) );
  INV_X1 U435 ( .A(KEYINPUT108), .ZN(n378) );
  NAND2_X1 U436 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U437 ( .A1(n381), .A2(n380), .ZN(n403) );
  INV_X1 U438 ( .A(n554), .ZN(n401) );
  XOR2_X1 U439 ( .A(KEYINPUT74), .B(G127GAT), .Z(n383) );
  XNOR2_X1 U440 ( .A(G78GAT), .B(G71GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U442 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n385) );
  XNOR2_X1 U443 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n399) );
  XOR2_X1 U446 ( .A(KEYINPUT73), .B(G64GAT), .Z(n389) );
  XNOR2_X1 U447 ( .A(G211GAT), .B(G183GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n394), .B(KEYINPUT76), .Z(n397) );
  XNOR2_X1 U453 ( .A(n395), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n580) );
  XOR2_X1 U456 ( .A(n580), .B(KEYINPUT107), .Z(n564) );
  INV_X1 U457 ( .A(n564), .ZN(n400) );
  NOR2_X1 U458 ( .A1(n401), .A2(n400), .ZN(n402) );
  AND2_X1 U459 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n404), .B(KEYINPUT47), .ZN(n411) );
  XOR2_X1 U461 ( .A(n554), .B(KEYINPUT95), .Z(n405) );
  XNOR2_X1 U462 ( .A(n405), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U463 ( .A1(n583), .A2(n580), .ZN(n406) );
  XNOR2_X1 U464 ( .A(KEYINPUT45), .B(n406), .ZN(n407) );
  NAND2_X1 U465 ( .A1(n407), .A2(n575), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n408), .B(KEYINPUT109), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n569), .B(KEYINPUT67), .ZN(n450) );
  INV_X1 U468 ( .A(n450), .ZN(n557) );
  NAND2_X1 U469 ( .A1(n409), .A2(n557), .ZN(n410) );
  NAND2_X1 U470 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n412), .B(KEYINPUT48), .ZN(n524) );
  XNOR2_X1 U472 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n413), .B(KEYINPUT85), .ZN(n414) );
  XOR2_X1 U474 ( .A(n414), .B(KEYINPUT21), .Z(n416) );
  XNOR2_X1 U475 ( .A(G197GAT), .B(G218GAT), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n432) );
  XNOR2_X1 U477 ( .A(n432), .B(n417), .ZN(n428) );
  XOR2_X1 U478 ( .A(n418), .B(G204GAT), .Z(n420) );
  NAND2_X1 U479 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT73), .Z(n422) );
  XNOR2_X1 U482 ( .A(G8GAT), .B(G169GAT), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U484 ( .A(n424), .B(n423), .Z(n426) );
  XNOR2_X1 U485 ( .A(G36GAT), .B(G92GAT), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n515) );
  NAND2_X1 U488 ( .A1(n524), .A2(n515), .ZN(n429) );
  XNOR2_X1 U489 ( .A(KEYINPUT54), .B(n429), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n443) );
  XOR2_X1 U491 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n434) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(G22GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(n435), .Z(n441) );
  XOR2_X1 U495 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n438) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U498 ( .A(KEYINPUT24), .B(n439), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n459) );
  NAND2_X1 U501 ( .A1(n568), .A2(n459), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U503 ( .A1(n527), .A2(n446), .ZN(n563) );
  NOR2_X1 U504 ( .A1(n554), .A2(n563), .ZN(n449) );
  XNOR2_X1 U505 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n471) );
  NAND2_X1 U506 ( .A1(n575), .A2(n450), .ZN(n485) );
  XOR2_X1 U507 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n452) );
  INV_X1 U508 ( .A(n580), .ZN(n479) );
  NAND2_X1 U509 ( .A1(n479), .A2(n554), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n468) );
  INV_X1 U511 ( .A(n518), .ZN(n529) );
  XOR2_X1 U512 ( .A(n515), .B(KEYINPUT27), .Z(n462) );
  NOR2_X1 U513 ( .A1(n462), .A2(n453), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n454), .B(KEYINPUT92), .ZN(n523) );
  NAND2_X1 U515 ( .A1(n529), .A2(n523), .ZN(n456) );
  XOR2_X1 U516 ( .A(n527), .B(KEYINPUT83), .Z(n455) );
  NOR2_X1 U517 ( .A1(n456), .A2(n455), .ZN(n467) );
  NAND2_X1 U518 ( .A1(n527), .A2(n515), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n459), .A2(n457), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n458), .B(KEYINPUT25), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n459), .A2(n527), .ZN(n460) );
  XNOR2_X1 U522 ( .A(KEYINPUT26), .B(n460), .ZN(n567) );
  INV_X1 U523 ( .A(n567), .ZN(n461) );
  NOR2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U525 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n513), .A2(n465), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n478) );
  NOR2_X1 U528 ( .A1(n468), .A2(n478), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT93), .ZN(n499) );
  NOR2_X1 U530 ( .A1(n485), .A2(n499), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n513), .A2(n476), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n515), .A2(n476), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT35), .B(KEYINPUT94), .Z(n474) );
  NAND2_X1 U536 ( .A1(n476), .A2(n527), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(n475), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n476), .A2(n518), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n477), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .Z(n488) );
  INV_X1 U542 ( .A(KEYINPUT97), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n479), .A2(n478), .ZN(n480) );
  XOR2_X1 U544 ( .A(KEYINPUT96), .B(n480), .Z(n481) );
  NOR2_X1 U545 ( .A1(n583), .A2(n481), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n484), .ZN(n512) );
  NOR2_X1 U548 ( .A1(n485), .A2(n512), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n486), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U550 ( .A1(n513), .A2(n495), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n495), .A2(n515), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n489), .B(KEYINPUT98), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n490), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n494) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n492) );
  NAND2_X1 U557 ( .A1(n527), .A2(n495), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT101), .Z(n497) );
  NAND2_X1 U561 ( .A1(n518), .A2(n495), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n502) );
  NAND2_X1 U564 ( .A1(n569), .A2(n375), .ZN(n511) );
  NOR2_X1 U565 ( .A1(n511), .A2(n499), .ZN(n500) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(n500), .Z(n508) );
  NAND2_X1 U567 ( .A1(n508), .A2(n513), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n505) );
  NAND2_X1 U571 ( .A1(n508), .A2(n515), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n508), .A2(n527), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U577 ( .A1(n508), .A2(n518), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n519) );
  NAND2_X1 U580 ( .A1(n513), .A2(n519), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n515), .A2(n519), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n527), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n522), .Z(G1339GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n545), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT111), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n532), .B(KEYINPUT113), .ZN(n533) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  NOR2_X1 U596 ( .A1(n542), .A2(n498), .ZN(n537) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n535) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n539) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  NOR2_X1 U604 ( .A1(n542), .A2(n564), .ZN(n540) );
  XOR2_X1 U605 ( .A(n541), .B(n540), .Z(G1342GAT) );
  NOR2_X1 U606 ( .A1(n542), .A2(n554), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n545), .A2(n567), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n569), .A2(n553), .ZN(n546) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n498), .A2(n553), .ZN(n551) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT52), .B(n549), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n580), .A2(n553), .ZN(n552) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT120), .B(n555), .Z(n556) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n563), .ZN(n558) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n498), .A2(n563), .ZN(n561) );
  XOR2_X1 U629 ( .A(n562), .B(n561), .Z(G1349GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n569), .A2(n582), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT124), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n582), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

