

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XOR2_X1 U326 ( .A(G57GAT), .B(KEYINPUT13), .Z(n369) );
  XNOR2_X1 U327 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U328 ( .A(n333), .B(n332), .Z(n514) );
  XOR2_X1 U329 ( .A(KEYINPUT21), .B(G211GAT), .Z(n294) );
  XOR2_X1 U330 ( .A(n370), .B(n328), .Z(n295) );
  OR2_X1 U331 ( .A1(n468), .A2(n572), .ZN(n296) );
  AND2_X1 U332 ( .A1(n465), .A2(n296), .ZN(n297) );
  XOR2_X1 U333 ( .A(G50GAT), .B(n496), .Z(n298) );
  XOR2_X1 U334 ( .A(KEYINPUT40), .B(n494), .Z(n299) );
  XNOR2_X1 U335 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n397) );
  XNOR2_X1 U336 ( .A(n398), .B(n397), .ZN(n570) );
  XNOR2_X1 U337 ( .A(n382), .B(n381), .ZN(n384) );
  XNOR2_X1 U338 ( .A(n439), .B(KEYINPUT55), .ZN(n454) );
  INV_X1 U339 ( .A(G190GAT), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n489), .B(KEYINPUT38), .ZN(n495) );
  XNOR2_X1 U341 ( .A(n455), .B(KEYINPUT58), .ZN(n456) );
  XNOR2_X1 U342 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n301) );
  XNOR2_X1 U344 ( .A(KEYINPUT9), .B(KEYINPUT79), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U346 ( .A(n302), .B(KEYINPUT66), .Z(n304) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n425) );
  XNOR2_X1 U348 ( .A(G134GAT), .B(n425), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n315) );
  XOR2_X1 U350 ( .A(KEYINPUT64), .B(KEYINPUT80), .Z(n306) );
  NAND2_X1 U351 ( .A1(G232GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U353 ( .A(n307), .B(KEYINPUT10), .Z(n313) );
  XOR2_X1 U354 ( .A(G29GAT), .B(G43GAT), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n356) );
  XOR2_X1 U357 ( .A(G92GAT), .B(G218GAT), .Z(n311) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n324) );
  XNOR2_X1 U360 ( .A(n356), .B(n324), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U363 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n317) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G85GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U366 ( .A(G99GAT), .B(n318), .ZN(n383) );
  XNOR2_X1 U367 ( .A(n319), .B(n383), .ZN(n388) );
  INV_X1 U368 ( .A(n388), .ZN(n555) );
  XNOR2_X1 U369 ( .A(n555), .B(KEYINPUT81), .ZN(n539) );
  XOR2_X1 U370 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n321) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n441) );
  XOR2_X1 U373 ( .A(G176GAT), .B(G64GAT), .Z(n370) );
  XOR2_X1 U374 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n327) );
  XNOR2_X1 U375 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n294), .B(n322), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n323), .B(G197GAT), .ZN(n436) );
  INV_X1 U378 ( .A(n436), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  NAND2_X1 U381 ( .A1(G226GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n295), .B(n329), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n441), .B(n330), .ZN(n333) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G183GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n331), .B(KEYINPUT82), .ZN(n340) );
  INV_X1 U386 ( .A(n340), .ZN(n332) );
  INV_X1 U387 ( .A(n514), .ZN(n461) );
  XOR2_X1 U388 ( .A(KEYINPUT84), .B(G64GAT), .Z(n335) );
  XNOR2_X1 U389 ( .A(G127GAT), .B(G71GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U391 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n337) );
  XNOR2_X1 U392 ( .A(KEYINPUT85), .B(KEYINPUT14), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n349) );
  XOR2_X1 U395 ( .A(G15GAT), .B(G1GAT), .Z(n353) );
  XOR2_X1 U396 ( .A(n340), .B(KEYINPUT83), .Z(n342) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n353), .B(n343), .ZN(n347) );
  XOR2_X1 U400 ( .A(n369), .B(G78GAT), .Z(n345) );
  XOR2_X1 U401 ( .A(G22GAT), .B(G155GAT), .Z(n422) );
  XNOR2_X1 U402 ( .A(G211GAT), .B(n422), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n583) );
  XOR2_X1 U406 ( .A(G22GAT), .B(G197GAT), .Z(n351) );
  XNOR2_X1 U407 ( .A(G50GAT), .B(G36GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U409 ( .A(n352), .B(G141GAT), .Z(n355) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(n353), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U412 ( .A(n356), .B(KEYINPUT70), .Z(n358) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U415 ( .A(n360), .B(n359), .Z(n368) );
  XOR2_X1 U416 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n362) );
  XNOR2_X1 U417 ( .A(G113GAT), .B(G8GAT), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n364) );
  XNOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n575) );
  XOR2_X1 U424 ( .A(n369), .B(G92GAT), .Z(n372) );
  XNOR2_X1 U425 ( .A(G204GAT), .B(n370), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U427 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n374) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n382) );
  XOR2_X1 U431 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  XOR2_X1 U432 ( .A(G148GAT), .B(G78GAT), .Z(n421) );
  XNOR2_X1 U433 ( .A(n440), .B(n421), .ZN(n380) );
  XOR2_X1 U434 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n378) );
  XNOR2_X1 U435 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n579) );
  XNOR2_X1 U438 ( .A(KEYINPUT41), .B(n579), .ZN(n564) );
  NOR2_X1 U439 ( .A1(n575), .A2(n564), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  NOR2_X1 U441 ( .A1(n583), .A2(n386), .ZN(n387) );
  NAND2_X1 U442 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n389), .B(KEYINPUT113), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT47), .ZN(n395) );
  XNOR2_X1 U445 ( .A(KEYINPUT36), .B(n539), .ZN(n587) );
  INV_X1 U446 ( .A(n583), .ZN(n568) );
  NOR2_X1 U447 ( .A1(n587), .A2(n568), .ZN(n391) );
  XOR2_X1 U448 ( .A(KEYINPUT45), .B(n391), .Z(n392) );
  NOR2_X1 U449 ( .A1(n579), .A2(n392), .ZN(n393) );
  NAND2_X1 U450 ( .A1(n393), .A2(n575), .ZN(n394) );
  NAND2_X1 U451 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U452 ( .A(KEYINPUT48), .B(n396), .ZN(n526) );
  NAND2_X1 U453 ( .A1(n461), .A2(n526), .ZN(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n400) );
  XNOR2_X1 U455 ( .A(G120GAT), .B(G148GAT), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U457 ( .A(G57GAT), .B(KEYINPUT4), .Z(n402) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U460 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U461 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n406) );
  NAND2_X1 U462 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(KEYINPUT5), .B(n407), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(G162GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U469 ( .A(n413), .B(n412), .Z(n420) );
  XOR2_X1 U470 ( .A(KEYINPUT0), .B(G134GAT), .Z(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT86), .B(G127GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U473 ( .A(G113GAT), .B(n416), .Z(n451) );
  XOR2_X1 U474 ( .A(KEYINPUT3), .B(KEYINPUT90), .Z(n418) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n429) );
  XNOR2_X1 U477 ( .A(n451), .B(n429), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n571) );
  INV_X1 U479 ( .A(n571), .ZN(n512) );
  XOR2_X1 U480 ( .A(G106GAT), .B(G218GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n435) );
  XOR2_X1 U484 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n428) );
  XNOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n433) );
  XOR2_X1 U487 ( .A(KEYINPUT88), .B(n429), .Z(n431) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n466) );
  NAND2_X1 U493 ( .A1(n512), .A2(n466), .ZN(n438) );
  OR2_X1 U494 ( .A1(n570), .A2(n438), .ZN(n439) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT20), .Z(n445) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U502 ( .A(G183GAT), .B(G190GAT), .Z(n449) );
  XNOR2_X1 U503 ( .A(G43GAT), .B(G99GAT), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n529) );
  NAND2_X1 U507 ( .A1(n454), .A2(n529), .ZN(n567) );
  NOR2_X1 U508 ( .A1(n539), .A2(n567), .ZN(n457) );
  NAND2_X1 U509 ( .A1(n461), .A2(n529), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n458), .A2(n466), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(KEYINPUT97), .ZN(n462) );
  XNOR2_X1 U514 ( .A(n462), .B(n461), .ZN(n468) );
  XNOR2_X1 U515 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n464) );
  NOR2_X1 U516 ( .A1(n529), .A2(n466), .ZN(n463) );
  XOR2_X1 U517 ( .A(n464), .B(n463), .Z(n572) );
  NOR2_X1 U518 ( .A1(n571), .A2(n297), .ZN(n471) );
  XNOR2_X1 U519 ( .A(n466), .B(KEYINPUT67), .ZN(n467) );
  XNOR2_X1 U520 ( .A(n467), .B(KEYINPUT28), .ZN(n527) );
  INV_X1 U521 ( .A(n529), .ZN(n516) );
  NOR2_X1 U522 ( .A1(n512), .A2(n468), .ZN(n525) );
  NAND2_X1 U523 ( .A1(n516), .A2(n525), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n527), .A2(n469), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n485) );
  NAND2_X1 U526 ( .A1(n583), .A2(n539), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT16), .B(n472), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n485), .A2(n473), .ZN(n499) );
  NOR2_X1 U529 ( .A1(n579), .A2(n575), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n474), .B(KEYINPUT78), .ZN(n488) );
  NAND2_X1 U531 ( .A1(n499), .A2(n488), .ZN(n483) );
  NOR2_X1 U532 ( .A1(n512), .A2(n483), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT34), .B(n475), .Z(n476) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n514), .A2(n483), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT100), .B(n477), .Z(n478) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(n478), .ZN(G1325GAT) );
  NOR2_X1 U538 ( .A1(n483), .A2(n516), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n480) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n527), .ZN(n522) );
  NOR2_X1 U544 ( .A1(n522), .A2(n483), .ZN(n484) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n484), .Z(G1327GAT) );
  NOR2_X1 U546 ( .A1(n587), .A2(n485), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n568), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT37), .ZN(n511) );
  NAND2_X1 U549 ( .A1(n488), .A2(n511), .ZN(n489) );
  NOR2_X1 U550 ( .A1(n495), .A2(n512), .ZN(n491) );
  XNOR2_X1 U551 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NOR2_X1 U554 ( .A1(n514), .A2(n495), .ZN(n493) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U556 ( .A1(n495), .A2(n516), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n299), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n495), .A2(n522), .ZN(n496) );
  XNOR2_X1 U559 ( .A(KEYINPUT104), .B(n298), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n501) );
  INV_X1 U563 ( .A(n575), .ZN(n544) );
  NOR2_X1 U564 ( .A1(n564), .A2(n544), .ZN(n510) );
  NAND2_X1 U565 ( .A1(n510), .A2(n499), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n512), .A2(n506), .ZN(n500) );
  XOR2_X1 U567 ( .A(n501), .B(n500), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n514), .A2(n506), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n516), .A2(n506), .ZN(n504) );
  XOR2_X1 U572 ( .A(KEYINPUT108), .B(n504), .Z(n505) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n505), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n506), .ZN(n508) );
  XNOR2_X1 U575 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NAND2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n521) );
  NOR2_X1 U579 ( .A1(n512), .A2(n521), .ZN(n513) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n521), .ZN(n515) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n521), .ZN(n517) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(n517), .Z(n518) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n520) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U590 ( .A(n524), .B(n523), .Z(G1339GAT) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n543) );
  NOR2_X1 U593 ( .A1(n527), .A2(n543), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n530), .ZN(n540) );
  NOR2_X1 U596 ( .A1(n575), .A2(n540), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  XNOR2_X1 U598 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n564), .A2(n540), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(n535), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n540), .A2(n568), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n546) );
  NOR2_X1 U610 ( .A1(n572), .A2(n543), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n556), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n553) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .Z(n551) );
  INV_X1 U617 ( .A(n564), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n556), .A2(n549), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n583), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n558) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NOR2_X1 U627 ( .A1(n575), .A2(n567), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT125), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT126), .Z(n563) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U632 ( .A(n563), .B(n562), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n564), .A2(n567), .ZN(n565) );
  XOR2_X1 U634 ( .A(n566), .B(n565), .Z(G1349GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n574) );
  INV_X1 U638 ( .A(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n575), .A2(n586), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n581) );
  INV_X1 U645 ( .A(n586), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n584), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

