//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(G116), .B(G119), .Z(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G116), .B(G119), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n196), .B2(new_n197), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n191), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT67), .B1(new_n189), .B2(new_n190), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n191), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT84), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT3), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G107), .ZN(new_n217));
  OR3_X1    g031(.A1(new_n209), .A2(KEYINPUT3), .A3(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(G101), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n215), .A2(new_n217), .A3(new_n223), .A4(new_n218), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n208), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n192), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n189), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n214), .B1(G104), .B2(new_n213), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n224), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n224), .B2(new_n233), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n205), .B(new_n231), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(G110), .B(G122), .Z(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n226), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n238), .A2(new_n244), .A3(new_n239), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G146), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT64), .A3(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(G146), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n247), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G125), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n249), .A2(G143), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(new_n251), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n254), .A3(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT0), .B(G128), .Z(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n252), .A2(new_n262), .A3(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n261), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT89), .B(G224), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n269), .B(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n243), .A2(new_n245), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n239), .B(KEYINPUT8), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n230), .A2(new_n276), .B1(KEYINPUT5), .B2(new_n197), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n276), .B2(new_n230), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n205), .B(new_n278), .C1(new_n235), .C2(new_n236), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n205), .A2(new_n231), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n224), .A2(new_n233), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n275), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT7), .B1(new_n271), .B2(G953), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n286));
  INV_X1    g100(.A(new_n261), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(G125), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n261), .A2(KEYINPUT91), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n269), .A2(new_n284), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n283), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n293), .B2(new_n242), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n274), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n274), .A2(new_n294), .A3(new_n296), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n188), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT9), .B(G234), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n260), .A2(new_n256), .ZN(new_n304));
  OAI211_X1 g118(.A(KEYINPUT10), .B(new_n304), .C1(new_n235), .C2(new_n236), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n225), .A2(new_n268), .A3(new_n221), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G137), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .A3(G134), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(G137), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT66), .B(G131), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(new_n311), .A3(new_n312), .A4(new_n309), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n255), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n260), .B1(new_n259), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n224), .A3(new_n233), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n305), .A2(new_n306), .A3(new_n318), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT69), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G227), .ZN(new_n330));
  XOR2_X1   g144(.A(new_n330), .B(KEYINPUT83), .Z(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G140), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n235), .A2(new_n236), .A3(new_n304), .ZN(new_n337));
  INV_X1    g151(.A(new_n321), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n317), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT12), .B1(new_n317), .B2(KEYINPUT86), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI221_X1 g155(.A(new_n317), .B1(KEYINPUT86), .B2(KEYINPUT12), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n324), .A2(KEYINPUT88), .A3(new_n333), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n305), .A2(new_n323), .A3(new_n306), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n317), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n333), .B1(new_n347), .B2(new_n324), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G469), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT72), .B(G902), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G902), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n333), .B1(new_n343), .B2(new_n324), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n324), .A3(new_n333), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n324), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n341), .B2(new_n342), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT87), .B(new_n361), .C1(new_n365), .C2(new_n333), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n351), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n300), .B(new_n303), .C1(new_n358), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n325), .A2(G952), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(G237), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n329), .B(new_n353), .C1(G234), .C2(G237), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT21), .B(G898), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G128), .B(G143), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT99), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n308), .ZN(new_n379));
  INV_X1    g193(.A(G122), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G116), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT98), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n227), .A2(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n213), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(G107), .A3(new_n383), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(KEYINPUT14), .A3(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n382), .A2(KEYINPUT14), .A3(G107), .A4(new_n383), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n379), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n378), .A2(new_n308), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n247), .A2(G128), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(G134), .C1(KEYINPUT13), .C2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n385), .A3(new_n386), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n302), .A2(new_n397), .A3(G953), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n395), .A3(new_n398), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(KEYINPUT100), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT100), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n403), .A3(new_n399), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n353), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT15), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n405), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G475), .ZN(new_n410));
  INV_X1    g224(.A(G237), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n327), .A2(G953), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n325), .A2(KEYINPUT69), .ZN(new_n413));
  OAI211_X1 g227(.A(G214), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n247), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n329), .A2(G143), .A3(G214), .A4(new_n411), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n315), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n315), .A3(new_n416), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n423));
  INV_X1    g237(.A(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G125), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT16), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n427), .A2(new_n424), .A3(KEYINPUT76), .A4(G125), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n257), .A2(G140), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n426), .B(new_n428), .C1(new_n427), .C2(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n431), .A2(new_n249), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n249), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n418), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n422), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT18), .A2(G131), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n415), .A2(new_n416), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n415), .A2(KEYINPUT93), .A3(new_n416), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n437), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n430), .A2(G146), .ZN(new_n444));
  XNOR2_X1  g258(.A(G125), .B(G140), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n249), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT92), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n417), .A2(new_n443), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n442), .A2(KEYINPUT94), .A3(new_n451), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n436), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(new_n209), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT96), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n422), .A2(new_n434), .A3(new_n435), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n442), .A2(KEYINPUT94), .A3(new_n451), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT94), .B1(new_n442), .B2(new_n451), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n458), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT96), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI22_X1  g279(.A1(new_n459), .A2(new_n465), .B1(new_n458), .B2(new_n456), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n410), .B1(new_n466), .B2(new_n355), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n454), .A2(new_n455), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n433), .B(KEYINPUT78), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n419), .A2(new_n421), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n445), .B1(KEYINPUT95), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n445), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n469), .B(new_n470), .C1(G146), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n458), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n459), .B2(new_n465), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT20), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n458), .B1(new_n468), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n463), .A2(new_n464), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n468), .A2(KEYINPUT96), .A3(new_n458), .A4(new_n460), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n485), .A2(G475), .A3(G902), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(new_n410), .A3(new_n355), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n485), .B2(KEYINPUT97), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n467), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n369), .A2(new_n375), .A3(new_n409), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n317), .A2(new_n265), .A3(new_n266), .A4(new_n267), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n310), .A2(G134), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n312), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n304), .A2(new_n316), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n500), .A3(KEYINPUT30), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n208), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n329), .A2(G210), .A3(new_n411), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(G101), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n202), .A2(new_n496), .A3(new_n207), .A4(new_n500), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT31), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n505), .A2(new_n513), .A3(new_n509), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n510), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n510), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n207), .A2(new_n202), .B1(new_n496), .B2(new_n500), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n509), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n495), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n519), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(KEYINPUT71), .A3(new_n512), .A4(new_n514), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n494), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n523), .A2(new_n526), .A3(new_n509), .A4(new_n527), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n353), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT73), .B(new_n353), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n505), .A2(new_n510), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n529), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n544), .A3(new_n538), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G472), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n534), .A2(new_n535), .ZN(new_n548));
  INV_X1    g362(.A(new_n533), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n525), .B2(new_n531), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n536), .A2(new_n547), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n329), .A2(G221), .A3(G234), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT22), .B(G137), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G119), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT23), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n559), .B2(G128), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n563), .B2(new_n560), .ZN(new_n564));
  XNOR2_X1  g378(.A(G119), .B(G128), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  AOI22_X1  g380(.A1(new_n564), .A2(G110), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n432), .B2(new_n433), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n433), .B(new_n569), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n564), .A2(G110), .B1(new_n565), .B2(new_n566), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT77), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n571), .A2(new_n572), .B1(new_n249), .B2(new_n445), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n572), .B2(new_n571), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n558), .B(new_n568), .C1(new_n570), .C2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n568), .B1(new_n574), .B2(new_n570), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n557), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n577), .A3(new_n353), .ZN(new_n578));
  NOR2_X1   g392(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n397), .B1(new_n353), .B2(G234), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT75), .Z(new_n583));
  NAND4_X1  g397(.A1(new_n575), .A2(new_n577), .A3(new_n353), .A4(new_n579), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n575), .A2(new_n577), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n582), .A2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT82), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n585), .A2(KEYINPUT82), .A3(new_n589), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n552), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n493), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n223), .ZN(G3));
  NAND2_X1  g411(.A1(new_n532), .A2(new_n353), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n352), .B1(new_n525), .B2(new_n531), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT101), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(G472), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT102), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n303), .B1(new_n358), .B2(new_n367), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n600), .A2(new_n607), .A3(G472), .A4(new_n602), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n604), .A2(new_n534), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n593), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT103), .Z(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n402), .A2(new_n612), .A3(new_n404), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n400), .A2(KEYINPUT33), .A3(new_n401), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n614), .A3(G478), .A4(new_n353), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n405), .A2(new_n406), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n487), .A2(new_n491), .ZN(new_n619));
  INV_X1    g433(.A(new_n467), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n300), .A2(new_n375), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n611), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT34), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NAND2_X1  g440(.A1(new_n488), .A2(new_n489), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n410), .A4(new_n355), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n620), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n409), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(KEYINPUT104), .A3(new_n375), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n620), .A2(new_n627), .A3(new_n630), .A4(new_n628), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n374), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n634), .A3(new_n300), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n611), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G107), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NAND4_X1  g452(.A1(new_n619), .A2(new_n375), .A3(new_n409), .A4(new_n620), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n368), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n534), .A3(new_n604), .A4(new_n608), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(KEYINPUT105), .ZN(new_n643));
  INV_X1    g457(.A(new_n576), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(KEYINPUT105), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n588), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n585), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT37), .B(G110), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT106), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n651), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n372), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(new_n371), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT107), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n633), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n552), .A2(new_n660), .A3(new_n369), .A4(new_n649), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XNOR2_X1  g476(.A(new_n658), .B(KEYINPUT39), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT40), .B1(new_n605), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n529), .B1(new_n521), .B2(new_n522), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n511), .A2(G472), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(G472), .A2(G902), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT108), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n536), .A2(new_n548), .A3(new_n551), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n298), .A2(new_n299), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT38), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n409), .A2(new_n188), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n492), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n665), .A2(new_n671), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n605), .A2(KEYINPUT40), .A3(new_n664), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n649), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n247), .ZN(G45));
  NOR3_X1   g494(.A1(new_n492), .A2(new_n618), .A3(new_n659), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n552), .A3(new_n369), .A4(new_n649), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NOR3_X1   g497(.A1(new_n492), .A2(new_n623), .A3(new_n618), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n324), .A2(KEYINPUT88), .A3(new_n333), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT88), .B1(new_n324), .B2(new_n333), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n348), .B1(new_n687), .B2(new_n343), .ZN(new_n688));
  OAI21_X1  g502(.A(G469), .B1(new_n688), .B2(new_n352), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n303), .A3(new_n354), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n689), .A2(new_n692), .A3(new_n303), .A4(new_n354), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n684), .A2(new_n552), .A3(new_n594), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND3_X1  g511(.A1(new_n552), .A2(new_n594), .A3(new_n694), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n635), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AND4_X1   g514(.A1(new_n375), .A2(new_n619), .A3(new_n409), .A4(new_n620), .ZN(new_n701));
  INV_X1    g515(.A(new_n672), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n690), .A2(new_n702), .A3(new_n188), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n701), .A2(new_n552), .A3(new_n649), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND2_X1  g519(.A1(new_n598), .A2(G472), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n533), .B1(new_n515), .B2(new_n524), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(KEYINPUT110), .A3(new_n590), .A4(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n590), .B(new_n707), .C1(new_n601), .C2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n374), .B1(new_n691), .B2(new_n693), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n492), .A2(new_n675), .A3(new_n702), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  AND2_X1   g531(.A1(new_n706), .A2(new_n707), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n681), .A2(new_n649), .A3(new_n703), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND3_X1  g534(.A1(new_n298), .A2(new_n187), .A3(new_n299), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n360), .A2(new_n362), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n354), .A3(new_n357), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(new_n303), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n621), .A2(new_n658), .A3(new_n722), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n548), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n547), .B1(new_n534), .B2(new_n535), .ZN(new_n729));
  OAI211_X1 g543(.A(KEYINPUT42), .B(new_n590), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT111), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n492), .A2(new_n618), .A3(new_n659), .A4(new_n721), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n585), .A2(new_n589), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n550), .A2(KEYINPUT32), .B1(new_n546), .B2(G472), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n548), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n736), .A3(new_n737), .A4(new_n726), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n725), .A2(new_n303), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n721), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n681), .A2(new_n552), .A3(new_n594), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n733), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  AND2_X1   g559(.A1(new_n552), .A2(new_n594), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n746), .A2(new_n660), .A3(new_n741), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n308), .ZN(G36));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n492), .A2(new_n749), .A3(new_n617), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n492), .B2(new_n617), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n604), .A2(new_n534), .A3(new_n608), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n649), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n722), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n363), .A2(new_n366), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(G469), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n357), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  INV_X1    g581(.A(new_n763), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(new_n356), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n763), .A2(KEYINPUT112), .A3(KEYINPUT46), .A4(new_n357), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n766), .A2(new_n769), .A3(new_n354), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n303), .A3(new_n663), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n755), .B2(new_n756), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT113), .B(new_n722), .C1(new_n755), .C2(new_n756), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n759), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n771), .A2(new_n777), .A3(new_n303), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n777), .B1(new_n771), .B2(new_n303), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n552), .A2(new_n594), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n732), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NAND3_X1  g597(.A1(new_n590), .A2(new_n303), .A3(new_n187), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n671), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n492), .A2(new_n617), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n689), .A2(new_n354), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT49), .Z(new_n790));
  OR4_X1    g604(.A1(new_n673), .A2(new_n787), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n747), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n620), .A2(new_n627), .A3(new_n628), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n409), .A2(new_n658), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n605), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n552), .A3(new_n649), .A4(new_n722), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n681), .A2(new_n649), .A3(new_n718), .A4(new_n741), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n744), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n704), .B1(new_n635), .B2(new_n698), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n695), .A2(new_n716), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n754), .A2(new_n493), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n596), .B1(new_n803), .B2(new_n649), .ZN(new_n804));
  INV_X1    g618(.A(new_n623), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n409), .B(new_n467), .C1(new_n487), .C2(new_n491), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n805), .B1(new_n621), .B2(new_n806), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n609), .A2(new_n593), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n799), .A2(new_n809), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n649), .A2(KEYINPUT115), .A3(new_n659), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT115), .B1(new_n649), .B2(new_n659), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n715), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n671), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n814), .A3(new_n740), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n682), .A2(new_n719), .A3(new_n661), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT52), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n682), .A2(new_n661), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n676), .A2(new_n672), .A3(new_n811), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n671), .A3(new_n726), .A4(new_n812), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n818), .A2(new_n820), .A3(new_n821), .A4(new_n719), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n810), .B2(new_n823), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n641), .A2(new_n650), .B1(new_n595), .B2(new_n493), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n609), .A2(new_n593), .A3(new_n807), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n747), .B1(new_n739), .B2(new_n743), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n802), .A4(new_n798), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n817), .A2(new_n822), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT54), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n690), .A2(new_n721), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n371), .A2(new_n834), .A3(new_n750), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n734), .B(new_n837), .C1(new_n548), .C2(new_n735), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT48), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n830), .B1(new_n829), .B2(new_n831), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT53), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n804), .A2(new_n808), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT116), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT116), .B1(new_n800), .B2(new_n801), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n823), .A3(new_n828), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n833), .A2(new_n839), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n838), .A2(KEYINPUT48), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n834), .A2(new_n371), .A3(new_n750), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n673), .A2(new_n187), .A3(new_n690), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n713), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n834), .A2(new_n713), .A3(new_n371), .A4(new_n750), .ZN(new_n857));
  INV_X1    g671(.A(new_n855), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT50), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n718), .A2(new_n649), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n853), .A2(new_n861), .A3(new_n835), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n671), .A2(new_n593), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n789), .A2(new_n303), .A3(new_n722), .A4(new_n371), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n671), .A2(new_n866), .A3(KEYINPUT118), .A4(new_n593), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n619), .A2(new_n620), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n617), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT120), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n753), .A2(new_n371), .A3(new_n713), .A4(new_n855), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n873), .A2(KEYINPUT50), .B1(new_n836), .B2(new_n861), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n865), .A2(new_n867), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(new_n864), .A3(new_n867), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n492), .A3(new_n618), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n878), .A3(new_n879), .A4(new_n856), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n303), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n789), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n778), .B2(new_n779), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT121), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n857), .A2(new_n721), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n887), .B(new_n883), .C1(new_n778), .C2(new_n779), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n852), .B1(new_n881), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT119), .B1(new_n863), .B2(new_n871), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n874), .A2(new_n878), .A3(new_n892), .A4(new_n856), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n895), .B(new_n896), .C1(new_n778), .C2(new_n779), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n886), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n894), .A2(new_n852), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n851), .B1(new_n890), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n876), .A2(new_n621), .A3(new_n877), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n853), .A2(new_n703), .A3(new_n713), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(G952), .A3(new_n325), .A4(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT122), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n850), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n791), .B1(new_n905), .B2(new_n906), .ZN(G75));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n840), .A2(new_n847), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n352), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n296), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n243), .A2(new_n245), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n273), .Z(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n913), .B(new_n914), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n329), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n915), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n908), .B(new_n919), .C1(new_n910), .C2(new_n296), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n918), .A3(new_n920), .ZN(G51));
  NAND2_X1  g735(.A1(new_n357), .A2(KEYINPUT57), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n357), .A2(KEYINPUT57), .ZN(new_n923));
  INV_X1    g737(.A(new_n849), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n848), .B1(new_n840), .B2(new_n847), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n350), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n909), .A2(new_n352), .A3(new_n768), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n917), .B1(new_n927), .B2(new_n928), .ZN(G54));
  NAND4_X1  g743(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .A4(new_n352), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n485), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n485), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n917), .ZN(G60));
  AND2_X1   g747(.A1(new_n613), .A2(new_n614), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n934), .B(new_n937), .C1(new_n924), .C2(new_n925), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n833), .B2(new_n849), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n938), .B(new_n918), .C1(new_n934), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(G63));
  NOR2_X1   g755(.A1(new_n646), .A2(new_n647), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n825), .A2(new_n826), .A3(new_n841), .ZN(new_n947));
  INV_X1    g761(.A(new_n801), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n699), .A3(new_n949), .A4(new_n704), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n947), .A2(new_n828), .A3(new_n846), .A4(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n831), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n943), .B(new_n946), .C1(new_n824), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n945), .B1(new_n840), .B2(new_n847), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n953), .B(new_n918), .C1(new_n587), .C2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n918), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n955), .A2(KEYINPUT61), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n917), .B1(new_n954), .B2(new_n943), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n909), .A2(new_n946), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n586), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n958), .B(new_n960), .C1(KEYINPUT124), .C2(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n957), .A2(new_n962), .ZN(G66));
  NAND2_X1  g777(.A1(new_n809), .A2(new_n329), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n271), .B2(new_n373), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n912), .B1(G898), .B2(new_n329), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  AND2_X1   g782(.A1(new_n503), .A2(new_n504), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(new_n474), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n715), .B(new_n590), .C1(new_n728), .C2(new_n729), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n772), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n828), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n816), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n775), .A2(new_n974), .A3(new_n782), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n971), .B1(new_n976), .B2(new_n329), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(G227), .B2(new_n329), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  OR3_X1    g793(.A1(new_n679), .A2(new_n816), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n679), .B2(new_n816), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n746), .B1(new_n621), .B2(new_n806), .ZN(new_n983));
  OR4_X1    g797(.A1(new_n605), .A2(new_n983), .A3(new_n664), .A4(new_n721), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n775), .A2(new_n982), .A3(new_n782), .A4(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n329), .A3(new_n971), .ZN(new_n986));
  INV_X1    g800(.A(G227), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n655), .B1(new_n971), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n978), .B(new_n986), .C1(new_n329), .C2(new_n988), .ZN(G72));
  XNOR2_X1  g803(.A(new_n668), .B(KEYINPUT63), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n976), .B2(new_n809), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  INV_X1    g807(.A(new_n543), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n991), .C1(new_n976), .C2(new_n809), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n993), .A2(new_n529), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n832), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n990), .B1(new_n998), .B2(new_n840), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n511), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n544), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n917), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n991), .B1(new_n985), .B2(new_n809), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n994), .A2(new_n529), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1005), .A2(KEYINPUT125), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT125), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1004), .A2(new_n1009), .ZN(G57));
endmodule


