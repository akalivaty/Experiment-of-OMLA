//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AND2_X1   g0007(.A1(G58), .A2(G232), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n208), .B(new_n212), .C1(G107), .C2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT66), .B(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n207), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n223), .A2(new_n228), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  AOI21_X1  g0049(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(G244), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G283), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n250), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  OAI211_X1 g0065(.A(G1), .B(G13), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT68), .A2(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT68), .A2(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(G45), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT5), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(G257), .B(new_n266), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT68), .A2(G1), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT68), .A2(G1), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT5), .B(G41), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n278), .A2(G274), .A3(new_n279), .A4(new_n266), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n263), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT83), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT83), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n263), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G200), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT84), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n252), .A2(new_n253), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT7), .B1(new_n289), .B2(new_n226), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n264), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(G107), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G77), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT6), .ZN(new_n299));
  INV_X1    g0099(.A(G97), .ZN(new_n300));
  INV_X1    g0100(.A(G107), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G97), .A2(G107), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(KEYINPUT6), .A3(G97), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n296), .B(new_n298), .C1(new_n226), .C2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n227), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n227), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(G13), .B(G20), .C1(new_n267), .C2(new_n268), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n276), .A2(new_n277), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G33), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G97), .ZN(new_n320));
  INV_X1    g0120(.A(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n300), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n283), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT84), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n284), .A2(new_n327), .A3(G200), .A4(new_n286), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n288), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n307), .A2(new_n309), .B1(new_n300), .B2(new_n321), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n283), .A2(G169), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n256), .A2(new_n258), .A3(new_n261), .A4(new_n260), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n281), .B1(new_n250), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G179), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n320), .A2(new_n330), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT78), .ZN(new_n338));
  INV_X1    g0138(.A(new_n314), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n226), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT72), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n215), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n226), .A2(new_n264), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n218), .A2(new_n226), .B1(new_n202), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n339), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT11), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT73), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n315), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n316), .A2(KEYINPUT73), .A3(G13), .A4(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n309), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n316), .A2(G20), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G68), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT12), .B1(new_n321), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n219), .A2(KEYINPUT12), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n347), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n257), .B1(G232), .B2(new_n251), .ZN(new_n363));
  NOR2_X1   g0163(.A1(G226), .A2(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n250), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n265), .A2(new_n275), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n316), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT76), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(new_n266), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n276), .A2(new_n277), .B1(new_n265), .B2(new_n275), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT76), .B1(new_n371), .B2(new_n250), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n372), .A3(G238), .ZN(new_n373));
  INV_X1    g0173(.A(G1), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n367), .A2(new_n374), .A3(G274), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT75), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n366), .A2(new_n373), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n361), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT14), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(KEYINPUT77), .A3(new_n380), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n377), .A2(KEYINPUT77), .A3(KEYINPUT13), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G179), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n360), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n359), .B1(new_n385), .B2(G190), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n378), .A2(new_n380), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G200), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n338), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(G169), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT14), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n381), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n359), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n388), .A2(new_n390), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(KEYINPUT78), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n351), .A2(new_n215), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT15), .B(G87), .Z(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n340), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT8), .B(G58), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n405), .A2(new_n344), .B1(new_n226), .B2(new_n215), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n309), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n352), .A2(new_n353), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n401), .B(new_n407), .C1(new_n408), .C2(new_n215), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n257), .A2(G232), .A3(new_n251), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n257), .A2(G238), .A3(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n301), .C2(new_n257), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n250), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n371), .A2(new_n250), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G244), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n375), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n409), .B1(G200), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n416), .A2(new_n324), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n392), .A2(new_n400), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT79), .ZN(new_n422));
  INV_X1    g0222(.A(G159), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n344), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n297), .A2(KEYINPUT79), .A3(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n201), .B1(new_n218), .B2(G58), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(new_n226), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n292), .A2(new_n226), .A3(new_n293), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT7), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n219), .B1(new_n431), .B2(new_n294), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n421), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G68), .B1(new_n290), .B2(new_n295), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n355), .A2(KEYINPUT66), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT66), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G68), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n437), .A3(G58), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n224), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(G20), .B1(new_n424), .B2(new_n425), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n434), .A2(new_n440), .A3(KEYINPUT16), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n433), .A2(new_n441), .A3(new_n309), .ZN(new_n442));
  INV_X1    g0242(.A(G58), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT8), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G58), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT71), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n445), .B2(G58), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n314), .B2(new_n353), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n446), .ZN(new_n451));
  INV_X1    g0251(.A(new_n444), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n321), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT80), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n315), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n312), .A2(new_n313), .B1(new_n316), .B2(G20), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n449), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G223), .A2(G1698), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n292), .B2(new_n293), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n251), .A2(G226), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n462), .A2(new_n463), .B1(G33), .B2(G87), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n464), .A2(new_n266), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n368), .A2(G232), .A3(new_n266), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(G190), .A3(new_n375), .A4(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n375), .C1(new_n464), .C2(new_n266), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G200), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n442), .A2(new_n460), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n442), .A2(new_n460), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n468), .A2(G169), .ZN(new_n478));
  INV_X1    g0278(.A(G179), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n468), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n477), .A2(KEYINPUT18), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT18), .B1(new_n477), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(new_n480), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT18), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n477), .A2(KEYINPUT18), .A3(new_n480), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n475), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n289), .A2(new_n215), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G222), .A2(G1698), .ZN(new_n492));
  XOR2_X1   g0292(.A(KEYINPUT69), .B(G223), .Z(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(G1698), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n250), .B(new_n491), .C1(new_n494), .C2(new_n289), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n414), .A2(G226), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n375), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n497), .A2(G179), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n203), .A2(G20), .ZN(new_n499));
  INV_X1    g0299(.A(G150), .ZN(new_n500));
  OAI221_X1 g0300(.A(new_n499), .B1(new_n500), .B2(new_n344), .C1(new_n342), .C2(new_n449), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n339), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n458), .A2(G50), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(new_n503), .C1(G50), .C2(new_n315), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n361), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n498), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT9), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n504), .A2(new_n507), .B1(G200), .B2(new_n497), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n495), .A2(G190), .A3(new_n496), .A4(new_n375), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT74), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT10), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT10), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n508), .A2(new_n509), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n506), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n416), .A2(G179), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n416), .A2(new_n361), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n409), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n490), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n420), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n301), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT23), .B1(new_n301), .B2(G20), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT87), .B1(new_n526), .B2(G20), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT87), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n528), .A2(new_n226), .A3(G33), .A4(G116), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(G20), .B1(new_n292), .B2(new_n293), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  OAI21_X1  g0333(.A(G87), .B1(new_n533), .B2(KEYINPUT86), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n532), .A2(new_n535), .B1(KEYINPUT86), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n226), .B1(new_n252), .B2(new_n253), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n537), .A2(new_n538), .A3(new_n534), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n531), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(KEYINPUT24), .B(new_n531), .C1(new_n536), .C2(new_n539), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n309), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n319), .A2(G107), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n315), .A2(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT25), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n250), .B1(new_n278), .B2(new_n279), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G264), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n550));
  OAI211_X1 g0350(.A(G250), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G294), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n250), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n554), .A3(new_n280), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n544), .A2(new_n545), .A3(new_n547), .A4(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n324), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT88), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n544), .A2(new_n562), .A3(new_n545), .A4(new_n547), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n555), .A2(G169), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n555), .A2(new_n479), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n559), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n278), .A2(G274), .A3(new_n266), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n269), .A2(G250), .A3(new_n266), .ZN(new_n571));
  INV_X1    g0371(.A(new_n526), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n292), .A2(new_n293), .B1(new_n216), .B2(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n220), .A2(new_n251), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n570), .B(new_n571), .C1(new_n575), .C2(new_n266), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n319), .A2(G87), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n226), .B1(new_n362), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n303), .A2(new_n210), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n340), .B2(new_n300), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n355), .C2(new_n537), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n403), .A2(new_n351), .B1(new_n584), .B2(new_n309), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n216), .A2(G1698), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n574), .B(new_n586), .C1(new_n252), .C2(new_n253), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n266), .B1(new_n587), .B2(new_n526), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(G190), .A3(new_n570), .A4(new_n571), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n577), .A2(new_n578), .A3(new_n585), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n351), .A2(new_n403), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n314), .A2(new_n315), .A3(new_n317), .A4(new_n402), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n584), .A2(new_n309), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n576), .A2(new_n361), .ZN(new_n596));
  INV_X1    g0396(.A(G274), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n269), .A2(new_n250), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n588), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n479), .A3(new_n571), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n591), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT85), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n591), .A2(new_n601), .A3(KEYINPUT85), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(G116), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n261), .B(new_n226), .C1(G33), .C2(new_n300), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(G20), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n309), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT20), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n608), .A2(KEYINPUT20), .A3(new_n309), .A4(new_n609), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n351), .A2(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n607), .B1(new_n316), .B2(G33), .ZN(new_n615));
  INV_X1    g0415(.A(new_n309), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n349), .A2(new_n615), .A3(new_n350), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n257), .A2(G257), .A3(new_n251), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n257), .A2(G264), .A3(G1698), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n289), .A2(G303), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n250), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n548), .A2(G270), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n280), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n618), .A2(G169), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n618), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(G200), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n623), .A2(G190), .A3(new_n280), .A4(new_n624), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n618), .A2(KEYINPUT21), .A3(G169), .A4(new_n625), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n623), .A2(new_n280), .A3(new_n624), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n618), .A3(G179), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n628), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n606), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n337), .A2(new_n522), .A3(new_n569), .A4(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n520), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n475), .B(new_n399), .C1(new_n387), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n486), .A2(new_n487), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n514), .A2(new_n516), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n506), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n522), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n602), .A2(KEYINPUT89), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n591), .A2(new_n601), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n557), .A2(new_n558), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n329), .A2(new_n649), .A3(new_n336), .A4(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n568), .A2(new_n560), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n628), .A2(new_n633), .A3(new_n635), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n263), .A2(new_n282), .A3(G179), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n361), .B1(new_n263), .B2(new_n282), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT90), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n331), .A2(new_n334), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n660), .A3(new_n323), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n649), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n604), .A2(new_n335), .A3(new_n605), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n666), .A3(new_n601), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n655), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n644), .B1(new_n645), .B2(new_n668), .ZN(G369));
  INV_X1    g0469(.A(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n316), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n652), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n564), .A2(new_n677), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n569), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n564), .A2(new_n568), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n653), .A2(new_n678), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT91), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n629), .A2(new_n678), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n653), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n636), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n688), .A2(new_n694), .ZN(G399));
  NOR2_X1   g0495(.A1(new_n581), .A2(G116), .ZN(new_n696));
  XOR2_X1   g0496(.A(new_n696), .B(KEYINPUT92), .Z(new_n697));
  INV_X1    g0497(.A(new_n229), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n697), .A2(new_n374), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n225), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n337), .A2(new_n569), .A3(new_n637), .A4(new_n678), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT31), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n599), .A2(new_n554), .A3(new_n549), .A4(new_n571), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n333), .B(G179), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n549), .A2(new_n554), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n710), .B2(new_n576), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n634), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT94), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n625), .B1(new_n708), .B2(new_n707), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT94), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n549), .A2(new_n554), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(KEYINPUT93), .A3(new_n571), .A4(new_n599), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n715), .A2(new_n716), .A3(new_n656), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n713), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n715), .A2(KEYINPUT30), .A3(new_n656), .A4(new_n718), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n634), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n283), .A3(new_n555), .A4(new_n576), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(new_n677), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n706), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n720), .A2(KEYINPUT95), .A3(new_n723), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT95), .B1(new_n720), .B2(new_n723), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT31), .B(new_n677), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n704), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n733), .B(new_n678), .C1(new_n655), .C2(new_n667), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n653), .B1(new_n564), .B2(new_n568), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n651), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n663), .B1(new_n662), .B2(new_n649), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n604), .A2(new_n663), .A3(new_n335), .A4(new_n605), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n601), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n677), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n734), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n703), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n374), .B1(new_n671), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n699), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT96), .B(G169), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n227), .B1(new_n749), .B2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n226), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n754), .A2(KEYINPUT98), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(KEYINPUT98), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n226), .A2(new_n324), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n479), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n757), .A2(G329), .B1(G322), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n752), .A2(new_n759), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n289), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(G303), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n226), .B1(new_n753), .B2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G294), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n479), .A2(new_n766), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n758), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n752), .A2(new_n767), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G326), .A2(new_n776), .B1(new_n778), .B2(G283), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n774), .A2(new_n752), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(KEYINPUT33), .A2(G317), .ZN(new_n782));
  AND2_X1   g0582(.A1(KEYINPUT33), .A2(G317), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n770), .A2(new_n773), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n768), .A2(new_n210), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G68), .B2(new_n781), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n778), .A2(G107), .ZN(new_n788));
  INV_X1    g0588(.A(new_n764), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G77), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n257), .B1(new_n760), .B2(new_n443), .C1(new_n202), .C2(new_n775), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT32), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n754), .B2(new_n423), .ZN(new_n794));
  INV_X1    g0594(.A(new_n754), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(KEYINPUT32), .A3(G159), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n792), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n791), .B(new_n797), .C1(new_n300), .C2(new_n771), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT97), .Z(new_n799));
  AOI21_X1  g0599(.A(new_n751), .B1(new_n785), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n750), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n698), .A2(new_n257), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n245), .B2(G45), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n701), .A2(new_n275), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(new_n808), .B1(new_n607), .B2(new_n698), .ZN(new_n809));
  NAND3_X1  g0609(.A1(G355), .A2(new_n229), .A3(new_n257), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n748), .B(new_n800), .C1(new_n804), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n803), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n691), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n692), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n747), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(G330), .B2(new_n691), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n520), .A2(new_n677), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n417), .A2(new_n418), .B1(new_n409), .B2(new_n677), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n639), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n678), .B(new_n824), .C1(new_n655), .C2(new_n667), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n668), .A2(new_n677), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n823), .B(KEYINPUT100), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(new_n732), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n748), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n748), .B1(new_n823), .B2(new_n801), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n750), .A2(new_n801), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G143), .A2(new_n761), .B1(new_n789), .B2(G159), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n835), .B2(new_n775), .C1(new_n500), .C2(new_n780), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n836), .A2(new_n837), .B1(G58), .B2(new_n772), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n757), .A2(G132), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n777), .A2(new_n355), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n289), .B(new_n841), .C1(G50), .C2(new_n769), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n257), .B1(new_n757), .B2(G311), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n776), .A2(G303), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G87), .A2(new_n778), .B1(new_n772), .B2(G97), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n301), .A2(new_n768), .B1(new_n780), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n760), .A2(new_n849), .B1(new_n764), .B2(new_n607), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n831), .B1(G77), .B2(new_n833), .C1(new_n751), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n830), .A2(new_n854), .ZN(G384));
  INV_X1    g0655(.A(KEYINPUT35), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n226), .B(new_n227), .C1(new_n306), .C2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n857), .B(G116), .C1(new_n856), .C2(new_n306), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT36), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n701), .A2(G77), .A3(new_n438), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(G50), .B2(new_n355), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n670), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n434), .A2(new_n440), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n314), .B1(new_n864), .B2(new_n421), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n441), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n456), .B1(new_n458), .B2(new_n449), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n675), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n450), .A2(new_n454), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n865), .B2(new_n441), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n872), .A2(KEYINPUT101), .A3(new_n675), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n489), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n477), .B1(new_n480), .B2(new_n869), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n470), .ZN(new_n878));
  INV_X1    g0678(.A(new_n480), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n470), .B1(new_n879), .B2(new_n872), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n870), .A2(new_n880), .A3(new_n873), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n881), .B2(new_n877), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n477), .A2(new_n869), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n475), .B2(new_n641), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n876), .A2(new_n470), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n877), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT40), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n359), .A2(new_n677), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n398), .A2(new_n399), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n387), .A2(new_n677), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n823), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n725), .B1(new_n705), .B2(KEYINPUT31), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT104), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n875), .B2(new_n882), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n897), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n727), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT104), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n900), .B1(new_n883), .B2(new_n889), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n895), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n899), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT105), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n522), .A2(new_n906), .ZN(new_n912));
  OAI21_X1  g0712(.A(G330), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT106), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n825), .A2(new_n821), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n397), .A2(new_n359), .B1(new_n390), .B2(new_n388), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n918), .A2(new_n892), .B1(new_n387), .B2(new_n677), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n921), .A2(new_n903), .B1(new_n641), .B2(new_n869), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n398), .A2(new_n677), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT39), .B1(new_n901), .B2(new_n902), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n883), .A2(new_n926), .A3(new_n889), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n642), .A2(new_n643), .ZN(new_n930));
  INV_X1    g0730(.A(new_n506), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n522), .B2(new_n742), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n929), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n935));
  XNOR2_X1  g0735(.A(new_n934), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n916), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n316), .A2(new_n671), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n859), .B1(new_n316), .B2(new_n862), .C1(new_n937), .C2(new_n938), .ZN(G367));
  NAND2_X1  g0739(.A1(new_n769), .A2(G116), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT46), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n940), .A2(new_n941), .B1(G311), .B2(new_n776), .ZN(new_n942));
  AOI22_X1  g0742(.A1(G303), .A2(new_n761), .B1(new_n789), .B2(G283), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n941), .C2(new_n940), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n780), .A2(new_n849), .B1(new_n777), .B2(new_n300), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n289), .B1(new_n771), .B2(new_n301), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(G317), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n948), .B2(new_n754), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n760), .A2(new_n500), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n771), .A2(new_n355), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n780), .A2(new_n423), .B1(new_n764), .B2(new_n202), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(G143), .C2(new_n776), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n289), .B1(new_n795), .B2(G137), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G58), .A2(new_n769), .B1(new_n778), .B2(G77), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n949), .B1(new_n950), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT112), .Z(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n750), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n578), .A2(new_n585), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n677), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n649), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n601), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n803), .A3(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n804), .B1(new_n229), .B2(new_n403), .C1(new_n240), .C2(new_n806), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT111), .Z(new_n967));
  NAND4_X1  g0767(.A1(new_n960), .A2(new_n965), .A3(new_n747), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n963), .A2(new_n964), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n323), .A2(new_n677), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n337), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT107), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n337), .A2(KEYINPUT107), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n661), .A2(new_n678), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n978), .B1(new_n975), .B2(new_n976), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n694), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n981), .B(new_n978), .C1(new_n975), .C2(new_n976), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n988), .A2(new_n989), .A3(new_n682), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n678), .B1(new_n990), .B2(new_n335), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n684), .A2(new_n686), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n980), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT42), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n999), .B(new_n986), .C1(new_n991), .C2(new_n995), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n971), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n982), .A2(new_n564), .A3(new_n568), .A4(new_n984), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n677), .B1(new_n1002), .B2(new_n336), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n993), .B(KEYINPUT42), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n997), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n986), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n996), .A2(new_n987), .A3(new_n997), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n970), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1001), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n687), .A2(new_n983), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n687), .A2(KEYINPUT44), .A3(new_n983), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1015));
  NAND3_X1  g0815(.A1(new_n688), .A2(new_n980), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1015), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n687), .B2(new_n983), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n693), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n684), .A2(new_n686), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT110), .B(new_n815), .C1(new_n1022), .C2(new_n992), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n681), .A2(new_n683), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n686), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n815), .A2(KEYINPUT110), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n815), .A2(KEYINPUT110), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1021), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n743), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1034), .A2(new_n694), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1020), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n743), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n699), .B(KEYINPUT41), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n746), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n968), .B1(new_n1009), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT113), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1038), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1036), .B2(new_n743), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1001), .B(new_n1008), .C1(new_n1044), .C2(new_n746), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1045), .A2(KEYINPUT113), .A3(new_n968), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1042), .A2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(new_n699), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1033), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1024), .A2(new_n813), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n697), .C1(G68), .C2(G77), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n405), .A2(G50), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT50), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n805), .B1(new_n237), .B2(new_n275), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n697), .A2(new_n229), .A3(new_n257), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1053), .A2(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n229), .A2(G107), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n804), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n289), .B1(new_n453), .B2(new_n781), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n423), .B2(new_n775), .C1(new_n403), .C2(new_n771), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n760), .A2(new_n202), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n355), .A2(new_n764), .B1(new_n777), .B2(new_n300), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n768), .A2(new_n215), .B1(new_n754), .B2(new_n500), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G322), .A2(new_n776), .B1(new_n781), .B2(G311), .ZN(new_n1067));
  INV_X1    g0867(.A(G303), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n764), .C1(new_n948), .C2(new_n760), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT48), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n847), .B2(new_n771), .C1(new_n849), .C2(new_n768), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT49), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n257), .B1(new_n795), .B2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n607), .B2(new_n777), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT114), .Z(new_n1075));
  AOI21_X1  g0875(.A(new_n1066), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n747), .B(new_n1060), .C1(new_n1076), .C2(new_n751), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1051), .B1(new_n745), .B2(new_n1031), .C1(new_n1052), .C2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n985), .A2(new_n803), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n804), .B1(new_n300), .B2(new_n229), .C1(new_n248), .C2(new_n806), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n775), .A2(new_n948), .B1(new_n760), .B2(new_n763), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT115), .Z(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n788), .B1(new_n849), .B2(new_n764), .C1(new_n1068), .C2(new_n780), .ZN(new_n1084));
  INV_X1    g0884(.A(G322), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1085), .A2(new_n754), .B1(new_n771), .B2(new_n607), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n257), .A3(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1083), .B(new_n1087), .C1(new_n847), .C2(new_n768), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT116), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n775), .A2(new_n500), .B1(new_n760), .B2(new_n423), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT51), .Z(new_n1091));
  NOR2_X1   g0891(.A1(new_n219), .A2(new_n768), .ZN(new_n1092));
  INV_X1    g0892(.A(G143), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n764), .A2(new_n405), .B1(new_n754), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n771), .A2(new_n215), .ZN(new_n1095));
  NOR4_X1   g0895(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n781), .A2(G50), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n257), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G87), .B2(new_n778), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n750), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1079), .A2(new_n747), .A3(new_n1080), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1020), .A2(new_n1035), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n745), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1048), .B1(new_n1102), .B2(new_n1050), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1036), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n875), .A2(new_n882), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n884), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n926), .B1(new_n1108), .B2(new_n883), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n927), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n748), .B1(new_n1111), .B2(new_n801), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n775), .A2(new_n847), .B1(new_n764), .B2(new_n300), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G107), .B2(new_n781), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT117), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n257), .B(new_n1115), .C1(G294), .C2(new_n757), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n607), .B2(new_n760), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1117), .A2(new_n786), .A3(new_n841), .A4(new_n1095), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n769), .A2(G150), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n289), .B1(new_n1119), .B2(KEYINPUT53), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT54), .B(G143), .Z(new_n1121));
  AOI22_X1  g0921(.A1(G128), .A2(new_n776), .B1(new_n789), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G132), .A2(new_n761), .B1(new_n778), .B2(G50), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n757), .A2(G125), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(KEYINPUT53), .B2(new_n1119), .C1(new_n423), .C2(new_n771), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G137), .C2(new_n781), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n750), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1112), .B(new_n1128), .C1(new_n453), .C2(new_n833), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n919), .B1(new_n825), .B2(new_n821), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n925), .B(new_n927), .C1(new_n1130), .C2(new_n923), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n731), .ZN(new_n1132));
  OAI211_X1 g0932(.A(G330), .B(new_n824), .C1(new_n1132), .C2(new_n896), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(new_n919), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n923), .B1(new_n883), .B2(new_n889), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n822), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n520), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n820), .B1(new_n741), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1138), .B2(new_n919), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1131), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n895), .B(G330), .C1(new_n896), .C2(new_n897), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1129), .B1(new_n1144), .B2(new_n745), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n522), .A2(new_n906), .A3(G330), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n742), .A2(new_n522), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n644), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n920), .B1(new_n732), .B2(new_n824), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n917), .B1(new_n1149), .B2(new_n1142), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n727), .A2(new_n731), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(G330), .A3(new_n824), .A4(new_n920), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n827), .C1(new_n896), .C2(new_n897), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n919), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1154), .A3(new_n1138), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1148), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1131), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1135), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n651), .A2(new_n735), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n661), .B1(new_n646), .B2(new_n648), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n601), .B(new_n738), .C1(new_n1160), .C2(new_n663), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n678), .B(new_n1137), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n919), .B1(new_n1162), .B2(new_n821), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n921), .A2(new_n924), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1111), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1157), .B1(new_n1166), .B2(new_n1142), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1048), .B1(new_n1156), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1148), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1152), .A2(new_n1154), .A3(new_n1138), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n917), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1133), .A2(new_n919), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n1141), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1169), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1144), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1145), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT120), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n933), .A2(new_n1179), .A3(new_n1146), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1148), .A2(KEYINPUT120), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1156), .B2(new_n1167), .ZN(new_n1183));
  AND4_X1   g0983(.A1(G330), .A2(new_n899), .A3(new_n904), .A4(new_n909), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n923), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n641), .A2(new_n869), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1108), .A2(new_n883), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1130), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n504), .A2(new_n869), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n517), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n517), .A2(new_n1189), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OR3_X1    g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT119), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1185), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1184), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1197), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n922), .B2(new_n928), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n899), .A2(new_n904), .A3(G330), .A4(new_n909), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1185), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1200), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1178), .B1(new_n1183), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1203), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1179), .B1(new_n933), .B2(new_n1146), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1179), .A2(new_n1146), .A3(new_n644), .A4(new_n1147), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1144), .B2(new_n1174), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n1214), .A3(KEYINPUT57), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1207), .A2(new_n1215), .A3(new_n699), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n833), .A2(G50), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n760), .A2(new_n301), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G41), .B(new_n257), .C1(new_n757), .C2(G283), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n778), .A2(G58), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n403), .C2(new_n764), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(G97), .C2(new_n781), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n951), .B1(G77), .B2(new_n769), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n607), .C2(new_n775), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT58), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n202), .B1(new_n252), .B2(G41), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G132), .A2(new_n781), .B1(new_n789), .B2(G137), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n776), .A2(G125), .B1(new_n772), .B2(G150), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n769), .A2(new_n1121), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n761), .A2(G128), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n778), .A2(G159), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G41), .B1(new_n795), .B2(G124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1233), .A2(new_n264), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1225), .B(new_n1226), .C1(new_n1232), .C2(new_n1236), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT118), .Z(new_n1238));
  AOI211_X1 g1038(.A(new_n748), .B(new_n1217), .C1(new_n1238), .C2(new_n750), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1194), .A2(new_n801), .A3(new_n1196), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1210), .A2(new_n746), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1216), .A2(new_n1241), .ZN(G375));
  NAND3_X1  g1042(.A1(new_n1150), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1174), .A2(new_n1243), .A3(new_n1038), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n757), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n289), .B1(new_n1245), .B2(new_n1068), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G107), .A2(new_n789), .B1(new_n772), .B2(new_n402), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n215), .B2(new_n777), .C1(new_n849), .C2(new_n775), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n760), .A2(new_n847), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n300), .A2(new_n768), .B1(new_n780), .B2(new_n607), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1246), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n757), .A2(G128), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n781), .A2(new_n1121), .B1(new_n772), .B2(G50), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n776), .A2(G132), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n257), .A3(new_n1220), .A4(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n760), .A2(new_n835), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n768), .A2(new_n423), .B1(new_n764), .B2(new_n500), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1252), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n750), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n747), .B(new_n1259), .C1(new_n920), .C2(new_n802), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n355), .B2(new_n832), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n746), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1244), .A2(new_n1263), .ZN(G381));
  AND3_X1   g1064(.A1(new_n1042), .A2(new_n1046), .A3(new_n1105), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G381), .A2(G384), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1268), .A2(KEYINPUT121), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1206), .B2(new_n745), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1048), .B1(new_n1272), .B2(new_n1178), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1271), .B1(new_n1273), .B2(new_n1215), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(KEYINPUT121), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1269), .A2(new_n1176), .A3(new_n1274), .A4(new_n1275), .ZN(G407));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1176), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(G343), .C2(new_n1277), .ZN(G409));
  XNOR2_X1  g1078(.A(G393), .B(G396), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1105), .B1(new_n1045), .B2(new_n968), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1265), .B2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1040), .A2(G390), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1282), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1176), .B1(new_n1216), .B2(new_n1241), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1210), .A2(new_n1214), .A3(new_n1038), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1241), .A2(new_n1176), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n676), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR4_X1   g1091(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1243), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1174), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT123), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1243), .A2(new_n1293), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(new_n1048), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT123), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(new_n1299), .A3(new_n1174), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1263), .ZN(new_n1302));
  INV_X1    g1102(.A(G384), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1301), .A2(G384), .A3(new_n1263), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1292), .A2(KEYINPUT125), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT125), .B1(new_n1292), .B2(new_n1306), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1241), .A2(new_n1176), .A3(new_n1287), .ZN(new_n1310));
  OAI211_X1 g1110(.A(KEYINPUT122), .B(new_n1310), .C1(new_n1274), .C2(new_n1176), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT122), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1306), .A2(new_n1311), .A3(new_n1313), .A4(new_n1290), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1289), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1285), .B1(new_n1309), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1291), .A2(G2897), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1317), .B(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G375), .A2(G378), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1290), .A3(new_n1310), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1320), .A2(KEYINPUT63), .A3(new_n1290), .A4(new_n1310), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1323), .B1(new_n1324), .B2(new_n1317), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1326), .B2(new_n1314), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1311), .A2(new_n1313), .A3(new_n1290), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT124), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1311), .A2(new_n1313), .A3(KEYINPUT124), .A4(new_n1290), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1319), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1327), .A2(new_n1332), .ZN(new_n1333));
  AOI22_X1  g1133(.A1(new_n1316), .A2(new_n1322), .B1(new_n1333), .B2(new_n1285), .ZN(G405));
  NAND3_X1  g1134(.A1(new_n1281), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1279), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1042), .A2(new_n1046), .A3(new_n1105), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1280), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1337), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1336), .B1(new_n1340), .B2(new_n1283), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1335), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT126), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1306), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1277), .A2(new_n1320), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1317), .A2(KEYINPUT126), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1345), .B1(new_n1344), .B2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1342), .A2(new_n1349), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1335), .B(new_n1341), .C1(new_n1348), .C2(new_n1346), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(G402));
endmodule


