//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G140), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT76), .ZN(new_n204));
  OR3_X1    g018(.A1(new_n202), .A2(KEYINPUT76), .A3(G125), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n199), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n198), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n207), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n202), .A2(KEYINPUT76), .A3(G125), .ZN(new_n210));
  XNOR2_X1  g024(.A(G125), .B(G140), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(KEYINPUT76), .ZN(new_n212));
  OAI211_X1 g026(.A(G146), .B(new_n209), .C1(new_n212), .C2(new_n199), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n197), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n218));
  OAI211_X1 g032(.A(G119), .B(new_n191), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n192), .B1(new_n215), .B2(new_n216), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n194), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G110), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n211), .B(KEYINPUT77), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n198), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n221), .A2(G110), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n195), .A2(new_n196), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n225), .B(new_n213), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT72), .B(G953), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT78), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT78), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n231), .A2(new_n234), .A3(G221), .A4(G234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n230), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n230), .A3(new_n235), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(G137), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n233), .A2(new_n230), .A3(new_n235), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(new_n236), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n229), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n223), .A2(new_n239), .A3(new_n228), .A4(new_n242), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n188), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n244), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n245), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n190), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n246), .A2(new_n189), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G116), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT69), .B1(new_n254), .B2(G119), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n193), .A3(G116), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n255), .B(new_n257), .C1(G116), .C2(new_n193), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT2), .B(G113), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n258), .B2(new_n259), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n258), .A2(new_n261), .A3(new_n259), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n198), .A2(G143), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G128), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT0), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n273));
  OR3_X1    g087(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n240), .A2(G134), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT65), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT11), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(G137), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n279), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(G134), .B(new_n240), .C1(new_n282), .C2(KEYINPUT11), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n278), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n279), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n289), .B(new_n291), .C1(new_n292), .C2(new_n286), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT68), .B1(new_n269), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT1), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n302), .A2(new_n272), .A3(new_n303), .A4(G128), .ZN(new_n304));
  INV_X1    g118(.A(new_n267), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n267), .A2(new_n268), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n191), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n297), .A2(new_n304), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n288), .A2(new_n278), .A3(new_n289), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n312));
  OAI211_X1 g126(.A(G131), .B(new_n311), .C1(new_n312), .C2(new_n286), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n295), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n295), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n265), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(KEYINPUT71), .B(new_n265), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(G101), .ZN(new_n324));
  INV_X1    g138(.A(G237), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n231), .A2(G210), .A3(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n324), .B(new_n326), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n264), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n329), .A2(new_n262), .B1(new_n259), .B2(new_n258), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n295), .A3(new_n314), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n322), .A2(KEYINPUT31), .A3(new_n328), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G472), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n320), .A2(new_n328), .A3(new_n331), .A4(new_n321), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT31), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n295), .A2(new_n314), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n295), .A2(new_n314), .A3(KEYINPUT73), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n330), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n265), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT28), .A3(new_n331), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n327), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n334), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n332), .A2(new_n333), .A3(new_n345), .A4(new_n188), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT32), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n349));
  AOI211_X1 g163(.A(new_n349), .B(new_n327), .C1(new_n341), .C2(new_n343), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n320), .A2(new_n331), .A3(new_n321), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n327), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n341), .A2(new_n343), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n353), .B2(new_n328), .ZN(new_n354));
  AOI211_X1 g168(.A(G902), .B(new_n350), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n348), .B1(new_n355), .B2(new_n333), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n354), .ZN(new_n357));
  INV_X1    g171(.A(new_n350), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n188), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT74), .A3(G472), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n253), .B1(new_n347), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G214), .B1(G237), .B2(G902), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT83), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G104), .ZN(new_n366));
  AND2_X1   g180(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n367));
  NOR2_X1   g181(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(G104), .A3(new_n365), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G101), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n369), .A2(new_n376), .A3(new_n371), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT81), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(KEYINPUT81), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT4), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n265), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n366), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT82), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n385), .B(G101), .C1(new_n387), .C2(new_n384), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n377), .A2(KEYINPUT81), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n329), .A2(new_n262), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n193), .A3(G116), .ZN(new_n394));
  OAI211_X1 g208(.A(G113), .B(new_n394), .C1(new_n258), .C2(new_n393), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(G110), .B(G122), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n383), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(new_n403), .A3(new_n398), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n277), .A2(G125), .ZN(new_n405));
  INV_X1    g219(.A(new_n309), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(G125), .ZN(new_n407));
  INV_X1    g221(.A(G953), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G224), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n402), .A2(new_n404), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(KEYINPUT7), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n407), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n392), .A2(new_n395), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n391), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n398), .B(KEYINPUT8), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n413), .B(new_n401), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n188), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G210), .B1(G237), .B2(G902), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT84), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n420), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n411), .A2(new_n188), .A3(new_n422), .A4(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n364), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(G234), .A2(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(G952), .A3(new_n408), .ZN(new_n426));
  INV_X1    g240(.A(new_n231), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(G902), .A3(new_n425), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT21), .B(G898), .Z(new_n429));
  OAI21_X1  g243(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n208), .A2(new_n213), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n433));
  AND2_X1   g247(.A1(KEYINPUT72), .A2(G953), .ZN(new_n434));
  NOR2_X1   g248(.A1(KEYINPUT72), .A2(G953), .ZN(new_n435));
  OAI211_X1 g249(.A(G214), .B(new_n325), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n266), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n231), .A2(G143), .A3(G214), .A4(new_n325), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND4_X1   g253(.A1(new_n433), .A2(new_n439), .A3(KEYINPUT17), .A4(G131), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n278), .B1(new_n437), .B2(new_n438), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n433), .B1(new_n441), .B2(KEYINPUT17), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n432), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n439), .B(G131), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n446), .A2(KEYINPUT17), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT88), .B(new_n432), .C1(new_n440), .C2(new_n442), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n372), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n204), .A2(new_n205), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n225), .B1(new_n198), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n441), .A2(new_n454), .A3(KEYINPUT18), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n454), .A2(KEYINPUT18), .A3(G131), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n453), .B(new_n455), .C1(new_n439), .C2(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n449), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n451), .B1(new_n449), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n188), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G475), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n451), .A3(new_n457), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n452), .A2(KEYINPUT19), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n224), .B2(KEYINPUT19), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n198), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n446), .B(new_n213), .C1(new_n465), .C2(KEYINPUT86), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(KEYINPUT86), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n457), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n451), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(KEYINPUT20), .A3(new_n472), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n461), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n478), .B2(G116), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(KEYINPUT89), .A2(G122), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT89), .A2(G122), .ZN(new_n483));
  OAI21_X1  g297(.A(G116), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n254), .A2(G122), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT90), .A3(KEYINPUT14), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n478), .A2(KEYINPUT14), .A3(G116), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n481), .A2(new_n484), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G107), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n365), .A3(new_n485), .ZN(new_n492));
  XNOR2_X1  g306(.A(G128), .B(G143), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n285), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(KEYINPUT91), .A3(G107), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n491), .A2(new_n492), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n484), .A2(new_n485), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G107), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n492), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n285), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(KEYINPUT13), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n266), .A2(G128), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(G134), .C1(KEYINPUT13), .C2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(KEYINPUT9), .A2(G234), .ZN(new_n506));
  NAND2_X1  g320(.A1(KEYINPUT9), .A2(G234), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT79), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT79), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n509), .A2(G217), .A3(new_n408), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n496), .A2(new_n504), .A3(new_n514), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n188), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT93), .ZN(new_n519));
  INV_X1    g333(.A(G478), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n516), .A2(new_n522), .A3(new_n188), .A4(new_n517), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n518), .A2(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n477), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n431), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G469), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n377), .B(KEYINPUT81), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n305), .A2(KEYINPUT1), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n297), .A2(new_n304), .A3(new_n308), .A4(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n388), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT10), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n381), .A2(new_n382), .A3(new_n277), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n290), .A2(new_n294), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n406), .A2(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n391), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n231), .A2(G227), .ZN(new_n542));
  XNOR2_X1  g356(.A(G110), .B(G140), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n534), .B1(new_n391), .B2(new_n309), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT12), .A3(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n531), .A2(new_n388), .A3(new_n533), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n309), .B1(new_n531), .B2(new_n388), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n545), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n547), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n544), .B1(new_n556), .B2(new_n541), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n530), .B(new_n188), .C1(new_n554), .C2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n546), .A2(KEYINPUT12), .A3(new_n547), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT12), .B1(new_n546), .B2(new_n547), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n541), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n544), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n545), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(G469), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(G469), .A2(G902), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n558), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n509), .A2(new_n188), .A3(new_n511), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n569), .A2(G221), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n362), .A2(new_n529), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  NOR2_X1   g389(.A1(new_n431), .A2(new_n572), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n332), .A2(new_n188), .A3(new_n345), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G472), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n346), .A3(new_n252), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT95), .B(G478), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n519), .A2(new_n523), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n517), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n514), .B1(new_n496), .B2(new_n504), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT33), .B1(new_n516), .B2(new_n517), .ZN(new_n586));
  OAI211_X1 g400(.A(G478), .B(new_n188), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n516), .A2(KEYINPUT33), .A3(new_n517), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n592), .A2(KEYINPUT94), .A3(G478), .A4(new_n188), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n581), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n579), .A2(new_n477), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT34), .B(G104), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  AOI21_X1  g411(.A(KEYINPUT20), .B1(new_n471), .B2(new_n472), .ZN(new_n598));
  INV_X1    g412(.A(new_n472), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n474), .B(new_n599), .C1(new_n462), .C2(new_n470), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n461), .A3(new_n526), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n579), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT35), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n239), .A2(new_n242), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(new_n229), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n229), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n188), .A4(new_n190), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n608), .A2(new_n229), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n229), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n188), .A3(new_n190), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n606), .B1(new_n618), .B2(new_n250), .ZN(new_n619));
  INV_X1    g433(.A(new_n250), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(KEYINPUT97), .A3(new_n617), .A4(new_n612), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n528), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n576), .A2(new_n623), .A3(new_n346), .A4(new_n578), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G110), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n624), .B(new_n626), .ZN(G12));
  INV_X1    g441(.A(KEYINPUT32), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n346), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n346), .A2(new_n628), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n352), .B2(new_n354), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n348), .B(new_n333), .C1(new_n631), .C2(new_n358), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT74), .B1(new_n359), .B2(G472), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n629), .B(new_n630), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n622), .A2(new_n572), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n426), .B(KEYINPUT99), .Z(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(G900), .B2(new_n428), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n602), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n634), .A2(new_n424), .A3(new_n635), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  NAND2_X1  g456(.A1(new_n351), .A2(new_n328), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n342), .A2(new_n327), .A3(new_n331), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n188), .ZN(new_n646));
  OAI21_X1  g460(.A(G472), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n347), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n638), .B(KEYINPUT39), .Z(new_n649));
  OAI21_X1  g463(.A(KEYINPUT40), .B1(new_n572), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n572), .A2(KEYINPUT40), .A3(new_n649), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n618), .A2(new_n250), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n364), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n421), .A2(new_n423), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n421), .A2(KEYINPUT38), .A3(new_n423), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n461), .A2(new_n475), .A3(new_n476), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n526), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n651), .A2(new_n655), .A3(new_n656), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NAND2_X1  g480(.A1(new_n589), .A2(new_n593), .ZN(new_n667));
  INV_X1    g481(.A(new_n581), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n662), .A2(new_n669), .A3(new_n638), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n634), .A2(new_n424), .A3(new_n635), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n657), .A2(new_n656), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n347), .B2(new_n361), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(KEYINPUT100), .A3(new_n635), .A4(new_n671), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  INV_X1    g493(.A(new_n431), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n594), .B1(new_n601), .B2(new_n461), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n530), .A2(KEYINPUT101), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n553), .A2(new_n548), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n564), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n541), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n534), .A2(new_n535), .B1(new_n539), .B2(new_n391), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n538), .B1(new_n687), .B2(new_n537), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n562), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n683), .B1(new_n690), .B2(new_n188), .ZN(new_n691));
  AOI211_X1 g505(.A(G902), .B(new_n682), .C1(new_n685), .C2(new_n689), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n692), .A3(new_n570), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n362), .A2(new_n680), .A3(new_n681), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT102), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  INV_X1    g511(.A(new_n602), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n362), .A2(new_n680), .A3(new_n698), .A4(new_n693), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NOR2_X1   g514(.A1(new_n554), .A2(new_n557), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n682), .B1(new_n701), .B2(G902), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n690), .A2(new_n188), .A3(new_n683), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n430), .A2(new_n702), .A3(new_n571), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n676), .A2(new_n623), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NOR3_X1   g520(.A1(new_n250), .A2(KEYINPUT103), .A3(new_n251), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT103), .B1(new_n250), .B2(new_n251), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n346), .A4(new_n578), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n578), .A2(new_n708), .A3(new_n346), .A4(new_n709), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n663), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(new_n704), .A3(new_n424), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n718), .B1(new_n715), .B2(new_n717), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n478), .ZN(G24));
  AND3_X1   g536(.A1(new_n578), .A2(new_n346), .A3(new_n654), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n702), .A2(new_n703), .A3(new_n571), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n675), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT106), .B1(new_n681), .B2(new_n638), .ZN(new_n726));
  AND4_X1   g540(.A1(KEYINPUT106), .A2(new_n662), .A3(new_n669), .A4(new_n638), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n723), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND3_X1  g543(.A1(new_n421), .A2(new_n656), .A3(new_n423), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT107), .B1(new_n572), .B2(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n421), .A2(new_n656), .A3(new_n423), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n571), .A4(new_n568), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n634), .A2(new_n252), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n670), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n681), .A2(KEYINPUT106), .A3(new_n638), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n629), .A2(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n629), .A2(KEYINPUT108), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n361), .A3(new_n630), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n710), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n731), .A4(new_n734), .ZN(new_n745));
  OAI22_X1  g559(.A1(new_n740), .A2(KEYINPUT42), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND4_X1  g561(.A1(new_n362), .A2(new_n640), .A3(new_n731), .A4(new_n734), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT109), .B(G134), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G36));
  AOI21_X1  g564(.A(new_n653), .B1(new_n578), .B2(new_n346), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT43), .B1(new_n477), .B2(new_n669), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n662), .A2(new_n753), .A3(new_n594), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT44), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n732), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT110), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n755), .A2(new_n761), .A3(new_n732), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT111), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n544), .B1(new_n684), .B2(new_n541), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n545), .A2(new_n688), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n563), .A2(KEYINPUT45), .A3(new_n565), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n769), .A3(G469), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n567), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n770), .B2(new_n567), .ZN(new_n772));
  INV_X1    g586(.A(new_n558), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n570), .A3(new_n649), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n757), .A2(new_n776), .A3(new_n760), .A4(new_n762), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n764), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  OAI22_X1  g593(.A1(new_n774), .A2(new_n570), .B1(KEYINPUT112), .B2(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n567), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n567), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n558), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n571), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n780), .A2(new_n671), .A3(new_n732), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n347), .A2(new_n361), .A3(new_n253), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n202), .ZN(G42));
  INV_X1    g606(.A(new_n754), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n753), .B1(new_n662), .B2(new_n594), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n637), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n724), .A2(new_n730), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n744), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT48), .Z(new_n799));
  AND2_X1   g613(.A1(new_n795), .A2(new_n715), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n780), .A2(new_n788), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n691), .A2(new_n692), .A3(new_n571), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n732), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n661), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT119), .B1(new_n693), .B2(new_n364), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n693), .A2(KEYINPUT119), .A3(new_n364), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n715), .A2(new_n806), .A3(new_n795), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  INV_X1    g623(.A(new_n797), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n808), .A2(new_n809), .B1(new_n723), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n806), .A2(new_n795), .A3(new_n715), .A4(new_n807), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT50), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n253), .A2(new_n426), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n796), .A2(new_n347), .A3(new_n647), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n477), .A3(new_n818), .A4(new_n594), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n803), .A2(new_n811), .A3(new_n813), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT121), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n809), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n723), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n813), .A2(new_n823), .A3(new_n824), .A4(new_n819), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT51), .A4(new_n803), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(new_n681), .A3(new_n818), .ZN(new_n829));
  INV_X1    g643(.A(G952), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n830), .B(G953), .C1(new_n820), .C2(new_n821), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n799), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n800), .A2(new_n725), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n675), .A2(new_n663), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n654), .A2(new_n639), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n648), .A2(new_n573), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(new_n641), .A3(new_n728), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n678), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n678), .A2(new_n837), .A3(KEYINPUT52), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n602), .B1(new_n681), .B2(KEYINPUT115), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(KEYINPUT115), .B2(new_n681), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n574), .B(new_n624), .C1(new_n579), .C2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n739), .A2(new_n723), .A3(new_n731), .A4(new_n734), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n748), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n634), .A2(new_n623), .A3(new_n638), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n572), .A3(new_n730), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n694), .A2(new_n699), .A3(new_n705), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n721), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n852), .A3(new_n746), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT53), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n641), .A2(new_n728), .A3(KEYINPUT116), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT116), .B1(new_n641), .B2(new_n728), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n678), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n840), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n746), .A3(new_n852), .A4(new_n850), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n860), .A3(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n852), .A2(new_n746), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n840), .B2(new_n858), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n852), .A2(new_n746), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n863), .A2(new_n865), .A3(new_n850), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n842), .B2(new_n853), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n832), .A2(new_n833), .A3(new_n861), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n830), .A2(new_n408), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n710), .A2(new_n656), .A3(new_n571), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n691), .A2(new_n692), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT49), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n477), .B(new_n669), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT113), .Z(new_n881));
  AOI21_X1  g695(.A(new_n648), .B1(new_n878), .B2(new_n877), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n661), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT114), .Z(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n884), .ZN(G75));
  NAND2_X1  g699(.A1(new_n868), .A2(new_n869), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G902), .A3(new_n420), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n402), .A2(new_n404), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n410), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT55), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n231), .A2(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G51));
  XOR2_X1   g709(.A(new_n567), .B(KEYINPUT57), .Z(new_n896));
  INV_X1    g710(.A(new_n872), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n871), .B1(new_n868), .B2(new_n869), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n690), .ZN(new_n900));
  INV_X1    g714(.A(new_n886), .ZN(new_n901));
  OR3_X1    g715(.A1(new_n901), .A2(new_n188), .A3(new_n770), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n894), .B1(new_n900), .B2(new_n902), .ZN(G54));
  NAND4_X1  g717(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n904));
  INV_X1    g718(.A(new_n471), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n894), .ZN(G60));
  OAI21_X1  g722(.A(new_n592), .B1(new_n897), .B2(new_n898), .ZN(new_n909));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n894), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n872), .B2(new_n861), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n592), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G63));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n917));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n868), .B2(new_n869), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n611), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n244), .A2(new_n245), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n913), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n917), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n920), .A2(new_n924), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(KEYINPUT61), .A3(new_n913), .A4(new_n921), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(G66));
  AOI21_X1  g743(.A(new_n408), .B1(new_n429), .B2(G224), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n721), .A2(new_n845), .A3(new_n851), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n932), .B2(new_n231), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n889), .B1(G898), .B2(new_n231), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  AOI21_X1  g750(.A(new_n231), .B1(G227), .B2(G900), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n316), .A2(new_n317), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(new_n464), .Z(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n427), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n362), .A2(new_n573), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n942), .A2(new_n844), .A3(new_n649), .A4(new_n730), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n791), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n678), .B(new_n665), .C1(new_n856), .C2(new_n857), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n641), .A2(new_n728), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT116), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n641), .A2(new_n728), .A3(KEYINPUT116), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n951), .A2(new_n952), .A3(new_n665), .A4(new_n678), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n778), .A2(new_n944), .A3(new_n946), .A4(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(KEYINPUT123), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(KEYINPUT123), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n941), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n775), .A2(new_n710), .A3(new_n834), .A4(new_n743), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT42), .B1(new_n735), .B2(new_n739), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n745), .A2(new_n744), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n958), .B(new_n748), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n678), .B1(new_n856), .B2(new_n857), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n791), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n427), .B1(new_n963), .B2(new_n778), .ZN(new_n964));
  INV_X1    g778(.A(new_n940), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n231), .A2(G900), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n938), .B1(new_n957), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n941), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n946), .A2(new_n953), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n778), .A4(new_n944), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n954), .A2(KEYINPUT123), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n967), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n937), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n957), .A2(new_n968), .A3(new_n938), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT124), .B1(new_n975), .B2(new_n967), .ZN(new_n979));
  INV_X1    g793(.A(new_n937), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n977), .A2(new_n981), .ZN(G72));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n963), .A2(new_n778), .A3(new_n931), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  AND3_X1   g800(.A1(new_n984), .A2(KEYINPUT125), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT125), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n322), .A2(new_n327), .A3(new_n331), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT126), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n987), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(new_n894), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n973), .A2(new_n974), .A3(new_n931), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n986), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n643), .A2(new_n854), .A3(new_n860), .A4(new_n989), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n995), .A2(new_n644), .B1(new_n986), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n988), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n984), .A2(KEYINPUT125), .A3(new_n986), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n999), .A3(new_n990), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(KEYINPUT127), .A3(new_n913), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n993), .A2(new_n997), .A3(new_n1001), .ZN(G57));
endmodule


