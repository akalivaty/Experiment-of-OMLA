//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n204));
  AND2_X1   g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G57gat), .A2(G64gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT93), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n203), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211));
  OAI221_X1 g010(.A(new_n202), .B1(new_n208), .B2(KEYINPUT93), .C1(new_n211), .C2(new_n204), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(G127gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(G155gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(G155gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n220), .B(KEYINPUT95), .Z(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n218), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G15gat), .ZN(new_n226));
  INV_X1    g025(.A(G22gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G15gat), .A2(G22gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT87), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT16), .B1(new_n228), .B2(new_n229), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(G1gat), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G1gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT16), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G8gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT88), .B(G8gat), .Z(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n241), .A3(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(KEYINPUT21), .B2(new_n213), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n224), .B1(new_n218), .B2(new_n219), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n225), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n225), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G99gat), .B(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT96), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G85gat), .A3(G92gat), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT7), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT7), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(KEYINPUT96), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT8), .ZN(new_n261));
  INV_X1    g060(.A(G85gat), .ZN(new_n262));
  INV_X1    g061(.A(G92gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n252), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT7), .ZN(new_n267));
  AOI22_X1  g066(.A1(KEYINPUT8), .A2(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n251), .A3(new_n259), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT97), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT14), .ZN(new_n272));
  INV_X1    g071(.A(G29gat), .ZN(new_n273));
  INV_X1    g072(.A(G36gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT84), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT83), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n279), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G29gat), .A2(G36gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n272), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n276), .A2(new_n278), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G29gat), .A2(G36gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT85), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n275), .A2(new_n277), .ZN(new_n287));
  XNOR2_X1  g086(.A(G43gat), .B(G50gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(KEYINPUT15), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n284), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(KEYINPUT15), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT17), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n290), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n285), .B(new_n297), .ZN(new_n298));
  OR3_X1    g097(.A1(new_n296), .A2(new_n289), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  NOR4_X1   g099(.A1(KEYINPUT84), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n282), .B1(new_n281), .B2(new_n272), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n278), .A2(new_n280), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G43gat), .B(G50gat), .Z(new_n306));
  INV_X1    g105(.A(KEYINPUT15), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n308), .A2(KEYINPUT86), .A3(new_n286), .A4(new_n287), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n292), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n296), .A2(new_n289), .A3(new_n298), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT17), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n271), .B1(new_n300), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT41), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n294), .A2(new_n299), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n266), .A2(new_n269), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G190gat), .B(G218gat), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OR4_X1    g121(.A1(KEYINPUT98), .A2(new_n313), .A3(new_n320), .A4(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n313), .B2(new_n320), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT17), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n295), .B1(new_n294), .B2(new_n299), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n321), .B(new_n319), .C1(new_n327), .C2(new_n271), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(KEYINPUT98), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n331));
  INV_X1    g130(.A(G134gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G162gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n324), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n338), .A3(new_n329), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n250), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G120gat), .B(G148gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G176gat), .B(G204gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G230gat), .A2(G233gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT101), .Z(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n269), .A2(KEYINPUT100), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n213), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n318), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n210), .A2(new_n212), .B1(new_n269), .B2(KEYINPUT100), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n270), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT10), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n214), .A2(new_n270), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n349), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n352), .A2(new_n348), .A3(new_n354), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n346), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT102), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT102), .B(new_n349), .C1(new_n355), .C2(new_n357), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT103), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n361), .A2(new_n346), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n343), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT66), .B(G183gat), .ZN(new_n374));
  INV_X1    g173(.A(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT67), .ZN(new_n377));
  NAND3_X1  g176(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n379), .A3(new_n382), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G169gat), .ZN(new_n387));
  INV_X1    g186(.A(G176gat), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT23), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT23), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n387), .A2(new_n388), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT25), .ZN(new_n394));
  INV_X1    g193(.A(new_n374), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT27), .ZN(new_n396));
  NOR2_X1   g195(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT28), .B(G190gat), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT27), .B(G183gat), .Z(new_n400));
  OAI21_X1  g199(.A(KEYINPUT28), .B1(new_n400), .B2(G190gat), .ZN(new_n401));
  NOR3_X1   g200(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n387), .B2(new_n388), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n401), .B(new_n381), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n383), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT64), .B1(new_n381), .B2(new_n382), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n378), .B1(G183gat), .B2(G190gat), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT25), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n411), .ZN(new_n412));
  OAI22_X1  g211(.A1(new_n399), .A2(new_n405), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n394), .A2(KEYINPUT68), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G113gat), .B(G120gat), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n416), .A2(KEYINPUT1), .ZN(new_n417));
  XNOR2_X1  g216(.A(G127gat), .B(G134gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT68), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n411), .B1(new_n386), .B2(new_n392), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n413), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n394), .A2(new_n414), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n421), .A3(new_n419), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT32), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n427), .B2(new_n428), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT69), .B(G15gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G43gat), .ZN(new_n433));
  XOR2_X1   g232(.A(G71gat), .B(G99gat), .Z(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  OAI221_X1 g236(.A(KEYINPUT32), .B1(new_n430), .B2(new_n437), .C1(new_n427), .C2(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n427), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT70), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n428), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n445), .A3(new_n428), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT71), .B1(new_n443), .B2(KEYINPUT34), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n439), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT29), .ZN(new_n450));
  XNOR2_X1  g249(.A(G155gat), .B(G162gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT2), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(G155gat), .B2(G162gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G141gat), .B(G148gat), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n452), .B(new_n451), .C1(new_n456), .C2(new_n455), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n450), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  XOR2_X1   g261(.A(G197gat), .B(G204gat), .Z(new_n463));
  AOI21_X1  g262(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G211gat), .B(G218gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT72), .B1(new_n463), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT72), .B(new_n466), .C1(new_n463), .C2(new_n464), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G228gat), .ZN(new_n473));
  INV_X1    g272(.A(G233gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n471), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT3), .B1(new_n476), .B2(new_n450), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n460), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n472), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT3), .B1(new_n467), .B2(new_n450), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n472), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G106gat), .ZN(new_n487));
  XOR2_X1   g286(.A(G50gat), .B(G78gat), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(KEYINPUT78), .B2(G22gat), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(G22gat), .B2(new_n489), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n485), .B(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n436), .A2(new_n438), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n443), .A2(KEYINPUT34), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n494), .A2(new_n497), .A3(new_n444), .A4(new_n446), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n449), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n420), .B(new_n478), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT3), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n419), .B1(new_n478), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n505), .B2(new_n478), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n478), .A2(new_n419), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n507), .B(new_n503), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n508), .B(KEYINPUT4), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(new_n503), .A3(new_n507), .A4(new_n512), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n504), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G1gat), .B(G29gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(new_n262), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT0), .B(G57gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  AND2_X1   g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n517), .B2(new_n521), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n517), .A2(KEYINPUT6), .A3(new_n521), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n425), .A2(G226gat), .A3(G233gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n422), .A2(new_n413), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(KEYINPUT29), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n471), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n531), .A3(new_n476), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G8gat), .B(G36gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G64gat), .B(G92gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT30), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541));
  INV_X1    g340(.A(new_n534), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n476), .B1(new_n528), .B2(new_n531), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n534), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n538), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n535), .B2(new_n538), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n499), .A2(new_n500), .A3(new_n527), .A4(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n527), .A2(new_n449), .A3(new_n493), .A4(new_n498), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT35), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n493), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT37), .ZN(new_n556));
  INV_X1    g355(.A(new_n538), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n543), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT79), .B(KEYINPUT37), .Z(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT38), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n525), .A2(new_n526), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT38), .B1(new_n535), .B2(KEYINPUT37), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n539), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n515), .A2(new_n507), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(G225gat), .A3(G233gat), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(KEYINPUT39), .ZN(new_n569));
  INV_X1    g368(.A(new_n521), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n501), .A2(new_n503), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(KEYINPUT39), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT40), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n522), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n549), .B(new_n575), .C1(new_n574), .C2(new_n573), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n555), .B1(new_n566), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n493), .A2(new_n563), .A3(new_n549), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n449), .A2(new_n498), .A3(KEYINPUT36), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT36), .B1(new_n449), .B2(new_n498), .ZN(new_n580));
  OAI22_X1  g379(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n554), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n243), .B1(new_n312), .B2(new_n300), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n317), .A2(new_n243), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT90), .B1(new_n588), .B2(KEYINPUT18), .ZN(new_n589));
  INV_X1    g388(.A(new_n243), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n325), .B2(new_n326), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(new_n586), .A3(new_n584), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n586), .A4(new_n584), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n600));
  INV_X1    g399(.A(G141gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT81), .B(G113gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n602), .B(new_n603), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n599), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n606), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n607), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n598), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT89), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n294), .A2(new_n240), .A3(new_n299), .A4(new_n242), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n584), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n586), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI211_X1 g420(.A(KEYINPUT89), .B(new_n619), .C1(new_n584), .C2(new_n617), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n597), .B(new_n615), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT91), .B1(new_n596), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n595), .A4(new_n589), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n592), .A2(new_n594), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n629), .B(new_n597), .C1(new_n621), .C2(new_n622), .ZN(new_n630));
  INV_X1    g429(.A(new_n615), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n582), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n582), .A2(KEYINPUT92), .A3(new_n633), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n373), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n563), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n549), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n549), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(G8gat), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n642), .B2(new_n646), .ZN(G1325gat));
  NAND2_X1  g446(.A1(new_n449), .A2(new_n498), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(G15gat), .B1(new_n638), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n579), .A2(new_n580), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n226), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n638), .B2(new_n653), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n555), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n582), .A2(new_n342), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT44), .ZN(new_n659));
  INV_X1    g458(.A(new_n342), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n554), .B2(new_n581), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n250), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n371), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n624), .A2(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n527), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n667), .A2(new_n660), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT104), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n636), .B2(new_n637), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n527), .A2(G29gat), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n674), .B2(new_n676), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(G1328gat));
  NOR2_X1   g478(.A1(new_n550), .A2(G36gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT105), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n670), .B2(new_n550), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(KEYINPUT46), .A3(new_n684), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(G1329gat));
  NOR2_X1   g489(.A1(new_n648), .A2(G43gat), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n674), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(G43gat), .ZN(new_n693));
  INV_X1    g492(.A(new_n669), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n659), .B2(new_n663), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n695), .B2(new_n651), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n692), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n692), .B2(new_n696), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1330gat));
  OAI21_X1  g499(.A(G50gat), .B1(new_n670), .B2(new_n493), .ZN(new_n701));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n674), .A2(new_n702), .A3(new_n555), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n701), .B2(new_n703), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(G1331gat));
  AND4_X1   g506(.A1(new_n668), .A2(new_n582), .A3(new_n343), .A4(new_n371), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n563), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g509(.A(new_n549), .B(KEYINPUT106), .Z(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(new_n716), .Z(G1333gat));
  NAND3_X1  g516(.A1(new_n708), .A2(G71gat), .A3(new_n651), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n649), .ZN(new_n719));
  INV_X1    g518(.A(G71gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n708), .B2(new_n649), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n555), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n633), .A2(new_n665), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n727), .B(KEYINPUT51), .C1(new_n661), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n582), .A2(new_n342), .A3(new_n728), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT110), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n730), .B2(new_n731), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n661), .A2(new_n735), .A3(KEYINPUT51), .A4(new_n728), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n563), .A2(new_n262), .A3(new_n371), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n668), .A2(new_n371), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n665), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n659), .B2(new_n663), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n563), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n738), .A2(new_n739), .B1(new_n262), .B2(new_n744), .ZN(G1336gat));
  NAND3_X1  g544(.A1(new_n711), .A2(new_n263), .A3(new_n371), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n737), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n263), .B1(new_n743), .B2(new_n549), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT52), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n664), .A2(new_n711), .A3(new_n741), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(new_n751), .B2(G92gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n746), .B1(new_n733), .B2(new_n737), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(KEYINPUT111), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755));
  AOI211_X1 g554(.A(new_n755), .B(new_n746), .C1(new_n733), .C2(new_n737), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n754), .B2(new_n756), .ZN(G1337gat));
  OR3_X1    g556(.A1(new_n648), .A2(G99gat), .A3(new_n372), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n651), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G99gat), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT112), .B1(new_n743), .B2(new_n651), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n738), .A2(new_n758), .B1(new_n760), .B2(new_n761), .ZN(G1338gat));
  INV_X1    g561(.A(G106gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n743), .B2(new_n555), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(KEYINPUT53), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n555), .A2(new_n763), .A3(new_n371), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT113), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n738), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n767), .B(KEYINPUT114), .Z(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n737), .B2(new_n747), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT53), .B1(new_n771), .B2(new_n764), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1339gat));
  NOR2_X1   g572(.A1(new_n618), .A2(new_n620), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT115), .Z(new_n775));
  AOI21_X1  g574(.A(new_n586), .B1(new_n591), .B2(new_n584), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n775), .A2(new_n776), .B1(new_n608), .B2(new_n610), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n628), .A2(new_n371), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n270), .A2(new_n213), .A3(new_n350), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n353), .A2(new_n270), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n356), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n357), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n348), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n364), .B2(new_n365), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n346), .B1(new_n358), .B2(KEYINPUT54), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n779), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n784), .A2(KEYINPUT54), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n783), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT102), .B1(new_n790), .B2(new_n349), .ZN(new_n791));
  INV_X1    g590(.A(new_n365), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n787), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n788), .B(new_n795), .C1(new_n370), .C2(new_n369), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n632), .B2(new_n628), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n660), .B1(new_n778), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n370), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n342), .A2(new_n801), .A3(new_n795), .A4(new_n788), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n628), .A2(new_n777), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n665), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n373), .A2(new_n633), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n806), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n802), .A2(new_n803), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n628), .A2(new_n371), .A3(new_n777), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n668), .B2(new_n796), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n660), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n808), .B(new_n809), .C1(new_n813), .C2(new_n665), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(new_n563), .A3(new_n499), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n712), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n633), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n371), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n665), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g622(.A1(new_n549), .A2(new_n660), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n816), .A2(new_n332), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n817), .A2(new_n342), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G134gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n827), .A2(new_n828), .A3(new_n830), .A4(new_n831), .ZN(G1343gat));
  NAND3_X1  g631(.A1(new_n807), .A2(new_n555), .A3(new_n814), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n651), .A2(new_n527), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n712), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n668), .A2(G141gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n786), .B2(new_n787), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n793), .A2(new_n843), .A3(new_n794), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n844), .A3(new_n779), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n633), .A2(new_n801), .A3(new_n845), .A4(new_n795), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n811), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n660), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n665), .B1(new_n848), .B2(new_n804), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n342), .B1(new_n846), .B2(new_n811), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n250), .B1(new_n852), .B2(new_n810), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n806), .B1(new_n853), .B2(KEYINPUT120), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n493), .A2(new_n840), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n841), .A2(KEYINPUT118), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n833), .A2(new_n858), .A3(new_n840), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n835), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n633), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n838), .B(new_n839), .C1(new_n861), .C2(new_n601), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n601), .B1(new_n860), .B2(new_n633), .ZN(new_n863));
  INV_X1    g662(.A(new_n838), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT58), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1344gat));
  XOR2_X1   g665(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n867));
  NAND2_X1  g666(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(new_n835), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n840), .B(new_n555), .C1(new_n849), .C2(new_n806), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n868), .A2(new_n371), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n867), .B1(new_n871), .B2(G148gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n841), .A2(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n856), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n859), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n371), .A3(new_n869), .ZN(new_n876));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n836), .A2(new_n877), .A3(new_n371), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  INV_X1    g682(.A(new_n878), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n860), .B2(new_n371), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n883), .B(new_n880), .C1(new_n885), .C2(new_n872), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n882), .A2(new_n886), .ZN(G1345gat));
  AOI21_X1  g686(.A(G155gat), .B1(new_n836), .B2(new_n665), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n665), .A2(G155gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n860), .B2(new_n889), .ZN(G1346gat));
  INV_X1    g689(.A(new_n833), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n891), .A2(new_n334), .A3(new_n824), .A4(new_n834), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n860), .A2(new_n342), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n334), .ZN(G1347gat));
  INV_X1    g693(.A(new_n552), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n815), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n549), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n668), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n711), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n633), .A2(new_n387), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT123), .ZN(G1348gat));
  NOR3_X1   g701(.A1(new_n897), .A2(new_n388), .A3(new_n372), .ZN(new_n903));
  INV_X1    g702(.A(new_n899), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n371), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n388), .B2(new_n905), .ZN(G1349gat));
  OR3_X1    g705(.A1(new_n899), .A2(new_n400), .A3(new_n250), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n395), .B1(new_n897), .B2(new_n250), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n904), .A2(new_n375), .A3(new_n342), .ZN(new_n914));
  OAI21_X1  g713(.A(G190gat), .B1(new_n897), .B2(new_n660), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT61), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(KEYINPUT61), .B2(new_n915), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n915), .B2(KEYINPUT61), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  AND2_X1   g719(.A1(new_n868), .A2(new_n870), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n652), .A2(new_n527), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n550), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n668), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n668), .A2(G197gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n922), .A2(new_n712), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n891), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT125), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n891), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n926), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n925), .A2(new_n934), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n372), .A2(G204gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n928), .A2(KEYINPUT62), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n371), .A3(new_n923), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G204gat), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT62), .B1(new_n928), .B2(new_n937), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .A4(new_n943), .ZN(G1353gat));
  OAI211_X1 g743(.A(new_n223), .B(new_n665), .C1(new_n930), .C2(new_n933), .ZN(new_n945));
  OAI21_X1  g744(.A(G211gat), .B1(new_n924), .B2(new_n250), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  AOI21_X1  g749(.A(new_n660), .B1(new_n929), .B2(new_n932), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n342), .A2(G218gat), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n951), .A2(G218gat), .B1(new_n924), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1355gat));
endmodule


