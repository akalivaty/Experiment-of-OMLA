

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708;

  BUF_X1 U362 ( .A(n528), .Z(n557) );
  XNOR2_X2 U363 ( .A(n535), .B(KEYINPUT19), .ZN(n518) );
  XNOR2_X2 U364 ( .A(n358), .B(G104), .ZN(n456) );
  XNOR2_X2 U365 ( .A(n414), .B(n413), .ZN(n682) );
  XNOR2_X2 U366 ( .A(n357), .B(n549), .ZN(n648) );
  NOR2_X1 U367 ( .A1(n706), .A2(n573), .ZN(n485) );
  INV_X1 U368 ( .A(n513), .ZN(n637) );
  INV_X2 U369 ( .A(G953), .ZN(n696) );
  NAND2_X1 U370 ( .A1(n610), .A2(n613), .ZN(n505) );
  NAND2_X1 U371 ( .A1(n528), .A2(n621), .ZN(n535) );
  INV_X2 U372 ( .A(n639), .ZN(n555) );
  INV_X1 U373 ( .A(G113), .ZN(n358) );
  NAND2_X2 U374 ( .A1(n350), .A2(n565), .ZN(n669) );
  AND2_X1 U375 ( .A1(n497), .A2(n496), .ZN(n499) );
  XNOR2_X1 U376 ( .A(n513), .B(n377), .ZN(n532) );
  XNOR2_X1 U377 ( .A(n387), .B(KEYINPUT71), .ZN(n421) );
  XNOR2_X1 U378 ( .A(n692), .B(G101), .ZN(n387) );
  BUF_X1 U379 ( .A(n692), .Z(n693) );
  XNOR2_X1 U380 ( .A(n445), .B(KEYINPUT4), .ZN(n692) );
  XNOR2_X2 U381 ( .A(n564), .B(KEYINPUT2), .ZN(n350) );
  XOR2_X1 U382 ( .A(KEYINPUT67), .B(G131), .Z(n458) );
  XNOR2_X1 U383 ( .A(n348), .B(G116), .ZN(n371) );
  INV_X1 U384 ( .A(G119), .ZN(n348) );
  INV_X1 U385 ( .A(KEYINPUT44), .ZN(n361) );
  XOR2_X1 U386 ( .A(G143), .B(G122), .Z(n457) );
  INV_X1 U387 ( .A(KEYINPUT79), .ZN(n347) );
  NAND2_X1 U388 ( .A1(n555), .A2(n492), .ZN(n487) );
  XOR2_X1 U389 ( .A(G137), .B(G113), .Z(n369) );
  XNOR2_X1 U390 ( .A(G128), .B(G119), .ZN(n400) );
  XOR2_X1 U391 ( .A(G107), .B(G104), .Z(n382) );
  NOR2_X1 U392 ( .A1(n545), .A2(n548), .ZN(n546) );
  NOR2_X1 U393 ( .A1(n544), .A2(n543), .ZN(n356) );
  XNOR2_X1 U394 ( .A(G137), .B(KEYINPUT68), .ZN(n691) );
  NOR2_X1 U395 ( .A1(n563), .A2(n562), .ZN(n695) );
  XNOR2_X1 U396 ( .A(n351), .B(KEYINPUT48), .ZN(n563) );
  XNOR2_X1 U397 ( .A(n359), .B(KEYINPUT45), .ZN(n675) );
  XNOR2_X1 U398 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U399 ( .A(n689), .B(n455), .ZN(n462) );
  OR2_X1 U400 ( .A1(n532), .A2(n487), .ZN(n411) );
  NAND2_X1 U401 ( .A1(n675), .A2(n695), .ZN(n564) );
  XNOR2_X1 U402 ( .A(n532), .B(n347), .ZN(n346) );
  NOR2_X1 U403 ( .A1(n513), .A2(n487), .ZN(n488) );
  XNOR2_X1 U404 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U405 ( .A(n520), .B(KEYINPUT111), .ZN(n521) );
  NOR2_X1 U406 ( .A1(n517), .A2(n516), .ZN(n550) );
  XNOR2_X1 U407 ( .A(n515), .B(n514), .ZN(n517) );
  XNOR2_X1 U408 ( .A(n375), .B(n374), .ZN(n567) );
  XNOR2_X1 U409 ( .A(n387), .B(n373), .ZN(n374) );
  XNOR2_X1 U410 ( .A(n402), .B(n362), .ZN(n403) );
  XNOR2_X1 U411 ( .A(n386), .B(n385), .ZN(n388) );
  XNOR2_X1 U412 ( .A(n384), .B(n383), .ZN(n385) );
  AND2_X1 U413 ( .A1(n343), .A2(n597), .ZN(n340) );
  XNOR2_X1 U414 ( .A(G110), .B(KEYINPUT16), .ZN(n341) );
  AND2_X1 U415 ( .A1(G214), .A2(n453), .ZN(n342) );
  XOR2_X1 U416 ( .A(KEYINPUT105), .B(n501), .Z(n343) );
  AND2_X1 U417 ( .A1(n431), .A2(n620), .ZN(n344) );
  XOR2_X1 U418 ( .A(n567), .B(KEYINPUT62), .Z(n345) );
  NAND2_X1 U419 ( .A1(n484), .A2(n470), .ZN(n574) );
  XNOR2_X2 U420 ( .A(n448), .B(n668), .ZN(n495) );
  NAND2_X1 U421 ( .A1(n632), .A2(n346), .ZN(n471) );
  XNOR2_X2 U422 ( .A(n376), .B(n566), .ZN(n513) );
  NAND2_X1 U423 ( .A1(n476), .A2(n493), .ZN(n477) );
  XNOR2_X2 U424 ( .A(n349), .B(n433), .ZN(n493) );
  NAND2_X1 U425 ( .A1(n518), .A2(n344), .ZN(n349) );
  XNOR2_X1 U426 ( .A(n350), .B(n619), .ZN(n659) );
  NAND2_X1 U427 ( .A1(n354), .A2(n352), .ZN(n351) );
  XNOR2_X1 U428 ( .A(n353), .B(KEYINPUT46), .ZN(n352) );
  NOR2_X2 U429 ( .A1(n707), .A2(n708), .ZN(n353) );
  XNOR2_X1 U430 ( .A(n356), .B(n355), .ZN(n354) );
  INV_X1 U431 ( .A(KEYINPUT69), .ZN(n355) );
  NAND2_X1 U432 ( .A1(n648), .A2(n550), .ZN(n551) );
  NOR2_X2 U433 ( .A1(n625), .A2(n624), .ZN(n357) );
  NAND2_X1 U434 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U435 ( .A1(n360), .A2(n340), .ZN(n359) );
  XNOR2_X1 U436 ( .A(n486), .B(n361), .ZN(n360) );
  BUF_X1 U437 ( .A(n592), .Z(n662) );
  XNOR2_X2 U438 ( .A(n499), .B(n498), .ZN(n613) );
  INV_X1 U439 ( .A(n669), .ZN(n592) );
  NOR2_X1 U440 ( .A1(n669), .A2(n575), .ZN(n579) );
  NOR2_X1 U441 ( .A1(n669), .A2(n566), .ZN(n568) );
  XNOR2_X1 U442 ( .A(n477), .B(KEYINPUT22), .ZN(n481) );
  XNOR2_X2 U443 ( .A(n367), .B(n366), .ZN(n445) );
  XOR2_X2 U444 ( .A(G122), .B(G107), .Z(n436) );
  XOR2_X1 U445 ( .A(n401), .B(n400), .Z(n362) );
  INV_X1 U446 ( .A(KEYINPUT72), .ZN(n506) );
  XNOR2_X1 U447 ( .A(n454), .B(n342), .ZN(n455) );
  NOR2_X1 U448 ( .A1(n475), .A2(n470), .ZN(n492) );
  XNOR2_X1 U449 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n396) );
  XNOR2_X1 U450 ( .A(KEYINPUT28), .B(KEYINPUT112), .ZN(n514) );
  NOR2_X1 U451 ( .A1(n524), .A2(n512), .ZN(n534) );
  XNOR2_X1 U452 ( .A(n462), .B(n461), .ZN(n577) );
  NOR2_X1 U453 ( .A1(G902), .A2(n577), .ZN(n463) );
  NOR2_X1 U454 ( .A1(n516), .A2(n640), .ZN(n525) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n593) );
  XOR2_X1 U456 ( .A(n464), .B(n463), .Z(n497) );
  XNOR2_X1 U457 ( .A(n490), .B(n489), .ZN(n612) );
  XNOR2_X1 U458 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U459 ( .A(G134), .B(n458), .ZN(n688) );
  XNOR2_X1 U460 ( .A(G146), .B(n688), .ZN(n378) );
  XOR2_X1 U461 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n364) );
  NOR2_X1 U462 ( .A1(G953), .A2(G237), .ZN(n453) );
  NAND2_X1 U463 ( .A1(n453), .A2(G210), .ZN(n363) );
  XNOR2_X1 U464 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U465 ( .A(n378), .B(n365), .ZN(n375) );
  XNOR2_X2 U466 ( .A(G143), .B(KEYINPUT64), .ZN(n367) );
  INV_X1 U467 ( .A(G128), .ZN(n366) );
  XNOR2_X1 U468 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n368) );
  XNOR2_X1 U469 ( .A(n369), .B(n368), .ZN(n372) );
  INV_X1 U470 ( .A(KEYINPUT3), .ZN(n370) );
  XNOR2_X1 U471 ( .A(n371), .B(n370), .ZN(n413) );
  XOR2_X1 U472 ( .A(n372), .B(n413), .Z(n373) );
  INV_X1 U473 ( .A(G902), .ZN(n447) );
  NAND2_X1 U474 ( .A1(n567), .A2(n447), .ZN(n376) );
  INV_X1 U475 ( .A(G472), .ZN(n566) );
  INV_X1 U476 ( .A(KEYINPUT6), .ZN(n377) );
  INV_X1 U477 ( .A(n378), .ZN(n386) );
  INV_X1 U478 ( .A(G110), .ZN(n379) );
  XNOR2_X1 U479 ( .A(n691), .B(n379), .ZN(n399) );
  XNOR2_X1 U480 ( .A(G140), .B(KEYINPUT76), .ZN(n380) );
  XNOR2_X1 U481 ( .A(n399), .B(n380), .ZN(n384) );
  NAND2_X1 U482 ( .A1(G227), .A2(n696), .ZN(n381) );
  XNOR2_X1 U483 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U484 ( .A(n388), .B(n421), .ZN(n664) );
  NOR2_X1 U485 ( .A1(G902), .A2(n664), .ZN(n390) );
  XNOR2_X1 U486 ( .A(KEYINPUT70), .B(G469), .ZN(n389) );
  XNOR2_X1 U487 ( .A(n390), .B(n389), .ZN(n491) );
  XNOR2_X1 U488 ( .A(n491), .B(KEYINPUT1), .ZN(n639) );
  XNOR2_X1 U489 ( .A(KEYINPUT15), .B(G902), .ZN(n423) );
  NAND2_X1 U490 ( .A1(G234), .A2(n423), .ZN(n391) );
  XNOR2_X1 U491 ( .A(KEYINPUT20), .B(n391), .ZN(n405) );
  NAND2_X1 U492 ( .A1(G221), .A2(n405), .ZN(n393) );
  XOR2_X1 U493 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n392) );
  XNOR2_X1 U494 ( .A(n393), .B(n392), .ZN(n634) );
  XNOR2_X1 U495 ( .A(n634), .B(KEYINPUT93), .ZN(n475) );
  INV_X1 U496 ( .A(G146), .ZN(n394) );
  XNOR2_X1 U497 ( .A(n394), .B(G125), .ZN(n418) );
  XNOR2_X1 U498 ( .A(n418), .B(G140), .ZN(n395) );
  XNOR2_X1 U499 ( .A(n395), .B(KEYINPUT10), .ZN(n689) );
  XNOR2_X1 U500 ( .A(n689), .B(n396), .ZN(n404) );
  NAND2_X1 U501 ( .A1(G234), .A2(n696), .ZN(n397) );
  XOR2_X1 U502 ( .A(KEYINPUT8), .B(n397), .Z(n442) );
  NAND2_X1 U503 ( .A1(G221), .A2(n442), .ZN(n398) );
  XNOR2_X1 U504 ( .A(n399), .B(n398), .ZN(n402) );
  XOR2_X1 U505 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n401) );
  NAND2_X1 U506 ( .A1(n593), .A2(n447), .ZN(n410) );
  NAND2_X1 U507 ( .A1(n405), .A2(G217), .ZN(n408) );
  XNOR2_X1 U508 ( .A(KEYINPUT25), .B(KEYINPUT91), .ZN(n406) );
  XNOR2_X1 U509 ( .A(n406), .B(KEYINPUT75), .ZN(n407) );
  XNOR2_X1 U510 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X2 U511 ( .A(n410), .B(n409), .ZN(n470) );
  XNOR2_X2 U512 ( .A(n411), .B(KEYINPUT33), .ZN(n630) );
  XNOR2_X1 U513 ( .A(n436), .B(n456), .ZN(n412) );
  XNOR2_X1 U514 ( .A(n412), .B(n341), .ZN(n414) );
  NAND2_X1 U515 ( .A1(n696), .A2(G224), .ZN(n415) );
  XNOR2_X1 U516 ( .A(n415), .B(KEYINPUT85), .ZN(n417) );
  XNOR2_X1 U517 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n416) );
  XNOR2_X1 U518 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U520 ( .A(n682), .B(n420), .ZN(n422) );
  XNOR2_X1 U521 ( .A(n422), .B(n421), .ZN(n585) );
  INV_X1 U522 ( .A(n423), .ZN(n565) );
  OR2_X2 U523 ( .A1(n585), .A2(n565), .ZN(n427) );
  INV_X1 U524 ( .A(G237), .ZN(n424) );
  NAND2_X1 U525 ( .A1(n447), .A2(n424), .ZN(n428) );
  NAND2_X1 U526 ( .A1(n428), .A2(G210), .ZN(n425) );
  XNOR2_X1 U527 ( .A(n425), .B(KEYINPUT87), .ZN(n426) );
  XNOR2_X2 U528 ( .A(n427), .B(n426), .ZN(n528) );
  NAND2_X1 U529 ( .A1(n428), .A2(G214), .ZN(n621) );
  XNOR2_X1 U530 ( .A(KEYINPUT88), .B(G898), .ZN(n677) );
  NOR2_X1 U531 ( .A1(n696), .A2(n677), .ZN(n685) );
  NAND2_X1 U532 ( .A1(n685), .A2(G902), .ZN(n429) );
  NAND2_X1 U533 ( .A1(n696), .A2(G952), .ZN(n509) );
  NAND2_X1 U534 ( .A1(n429), .A2(n509), .ZN(n431) );
  NAND2_X1 U535 ( .A1(G237), .A2(G234), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n430), .B(KEYINPUT14), .ZN(n620) );
  INV_X1 U537 ( .A(KEYINPUT84), .ZN(n432) );
  XNOR2_X1 U538 ( .A(n432), .B(KEYINPUT0), .ZN(n433) );
  NAND2_X1 U539 ( .A1(n630), .A2(n493), .ZN(n435) );
  INV_X1 U540 ( .A(KEYINPUT34), .ZN(n434) );
  XNOR2_X1 U541 ( .A(n435), .B(n434), .ZN(n467) );
  XNOR2_X1 U542 ( .A(G116), .B(n436), .ZN(n437) );
  XNOR2_X1 U543 ( .A(n437), .B(KEYINPUT103), .ZN(n441) );
  XOR2_X1 U544 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n439) );
  XNOR2_X1 U545 ( .A(G134), .B(KEYINPUT102), .ZN(n438) );
  XNOR2_X1 U546 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U547 ( .A(n441), .B(n440), .Z(n444) );
  NAND2_X1 U548 ( .A1(G217), .A2(n442), .ZN(n443) );
  XNOR2_X1 U549 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U550 ( .A(n446), .B(n445), .ZN(n670) );
  NAND2_X1 U551 ( .A1(n670), .A2(n447), .ZN(n448) );
  INV_X1 U552 ( .A(G478), .ZN(n668) );
  XOR2_X1 U553 ( .A(KEYINPUT13), .B(KEYINPUT100), .Z(n450) );
  XNOR2_X1 U554 ( .A(KEYINPUT101), .B(G475), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n450), .B(n449), .ZN(n464) );
  XOR2_X1 U556 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n452) );
  XNOR2_X1 U557 ( .A(KEYINPUT12), .B(KEYINPUT99), .ZN(n451) );
  XNOR2_X1 U558 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U559 ( .A(n456), .B(KEYINPUT98), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n458), .B(n457), .ZN(n459) );
  NOR2_X1 U561 ( .A1(n495), .A2(n497), .ZN(n465) );
  XOR2_X1 U562 ( .A(n465), .B(KEYINPUT108), .Z(n527) );
  XNOR2_X1 U563 ( .A(n527), .B(KEYINPUT77), .ZN(n466) );
  NAND2_X1 U564 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U565 ( .A(n468), .B(KEYINPUT35), .ZN(n706) );
  INV_X1 U566 ( .A(KEYINPUT86), .ZN(n469) );
  XNOR2_X1 U567 ( .A(n639), .B(n469), .ZN(n537) );
  INV_X1 U568 ( .A(n537), .ZN(n472) );
  XOR2_X1 U569 ( .A(KEYINPUT107), .B(n470), .Z(n632) );
  NOR2_X1 U570 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U571 ( .A(KEYINPUT78), .B(n473), .Z(n478) );
  NAND2_X1 U572 ( .A1(n497), .A2(n495), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n474), .B(KEYINPUT106), .ZN(n624) );
  NOR2_X1 U574 ( .A1(n624), .A2(n475), .ZN(n476) );
  NOR2_X1 U575 ( .A1(n478), .A2(n481), .ZN(n480) );
  XOR2_X1 U576 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n479) );
  XNOR2_X1 U577 ( .A(n480), .B(n479), .ZN(n573) );
  NOR2_X2 U578 ( .A1(n481), .A2(n555), .ZN(n504) );
  NAND2_X1 U579 ( .A1(n504), .A2(n513), .ZN(n482) );
  XNOR2_X1 U580 ( .A(KEYINPUT66), .B(n482), .ZN(n483) );
  INV_X1 U581 ( .A(n483), .ZN(n484) );
  NAND2_X1 U582 ( .A1(n485), .A2(n574), .ZN(n486) );
  XOR2_X1 U583 ( .A(KEYINPUT95), .B(n488), .Z(n646) );
  NAND2_X1 U584 ( .A1(n646), .A2(n493), .ZN(n490) );
  XOR2_X1 U585 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n489) );
  BUF_X1 U586 ( .A(n491), .Z(n516) );
  INV_X1 U587 ( .A(n492), .ZN(n640) );
  AND2_X1 U588 ( .A1(n525), .A2(n513), .ZN(n494) );
  NAND2_X1 U589 ( .A1(n494), .A2(n493), .ZN(n600) );
  NAND2_X1 U590 ( .A1(n612), .A2(n600), .ZN(n500) );
  INV_X1 U591 ( .A(n495), .ZN(n496) );
  OR2_X1 U592 ( .A1(n496), .A2(n497), .ZN(n610) );
  INV_X1 U593 ( .A(KEYINPUT104), .ZN(n498) );
  NAND2_X1 U594 ( .A1(n500), .A2(n505), .ZN(n501) );
  INV_X1 U595 ( .A(n532), .ZN(n502) );
  NOR2_X1 U596 ( .A1(n632), .A2(n502), .ZN(n503) );
  NAND2_X1 U597 ( .A1(n504), .A2(n503), .ZN(n597) );
  INV_X1 U598 ( .A(n505), .ZN(n626) );
  NOR2_X1 U599 ( .A1(KEYINPUT47), .A2(n626), .ZN(n507) );
  XNOR2_X1 U600 ( .A(n507), .B(n506), .ZN(n519) );
  NOR2_X1 U601 ( .A1(G900), .A2(n696), .ZN(n508) );
  NAND2_X1 U602 ( .A1(n508), .A2(G902), .ZN(n510) );
  NAND2_X1 U603 ( .A1(n510), .A2(n509), .ZN(n511) );
  NAND2_X1 U604 ( .A1(n511), .A2(n620), .ZN(n524) );
  NAND2_X1 U605 ( .A1(n634), .A2(n470), .ZN(n512) );
  NAND2_X1 U606 ( .A1(n534), .A2(n637), .ZN(n515) );
  NAND2_X1 U607 ( .A1(n550), .A2(n518), .ZN(n607) );
  NOR2_X1 U608 ( .A1(n519), .A2(n607), .ZN(n531) );
  NAND2_X1 U609 ( .A1(n637), .A2(n621), .ZN(n522) );
  XOR2_X1 U610 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n520) );
  NOR2_X1 U611 ( .A1(n524), .A2(n523), .ZN(n526) );
  NAND2_X1 U612 ( .A1(n526), .A2(n525), .ZN(n545) );
  OR2_X1 U613 ( .A1(n545), .A2(n527), .ZN(n530) );
  INV_X1 U614 ( .A(n557), .ZN(n529) );
  NOR2_X1 U615 ( .A1(n530), .A2(n529), .ZN(n572) );
  NOR2_X1 U616 ( .A1(n531), .A2(n572), .ZN(n539) );
  NOR2_X1 U617 ( .A1(n532), .A2(n610), .ZN(n533) );
  NAND2_X1 U618 ( .A1(n534), .A2(n533), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n552), .A2(n535), .ZN(n536) );
  XNOR2_X1 U620 ( .A(n536), .B(KEYINPUT36), .ZN(n538) );
  NAND2_X1 U621 ( .A1(n538), .A2(n537), .ZN(n617) );
  NAND2_X1 U622 ( .A1(n539), .A2(n617), .ZN(n544) );
  NAND2_X1 U623 ( .A1(n607), .A2(KEYINPUT47), .ZN(n540) );
  XNOR2_X1 U624 ( .A(n540), .B(KEYINPUT80), .ZN(n542) );
  NAND2_X1 U625 ( .A1(n626), .A2(KEYINPUT47), .ZN(n541) );
  NAND2_X1 U626 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U627 ( .A(n557), .B(KEYINPUT38), .ZN(n548) );
  XNOR2_X1 U628 ( .A(n546), .B(KEYINPUT39), .ZN(n560) );
  NOR2_X1 U629 ( .A1(n560), .A2(n610), .ZN(n547) );
  XNOR2_X1 U630 ( .A(n547), .B(KEYINPUT40), .ZN(n708) );
  INV_X1 U631 ( .A(n548), .ZN(n622) );
  XNOR2_X1 U632 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n549) );
  XOR2_X1 U633 ( .A(KEYINPUT42), .B(n551), .Z(n707) );
  INV_X1 U634 ( .A(n552), .ZN(n553) );
  NAND2_X1 U635 ( .A1(n553), .A2(n621), .ZN(n554) );
  NOR2_X1 U636 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U637 ( .A(n556), .B(KEYINPUT43), .ZN(n558) );
  NOR2_X1 U638 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U639 ( .A(n559), .B(KEYINPUT109), .ZN(n705) );
  NOR2_X1 U640 ( .A1(n613), .A2(n560), .ZN(n618) );
  INV_X1 U641 ( .A(n618), .ZN(n561) );
  NAND2_X1 U642 ( .A1(n705), .A2(n561), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n568), .B(n345), .ZN(n570) );
  INV_X1 U644 ( .A(G952), .ZN(n569) );
  AND2_X1 U645 ( .A1(n569), .A2(G953), .ZN(n674) );
  NAND2_X1 U646 ( .A1(n570), .A2(n588), .ZN(n571) );
  XNOR2_X1 U647 ( .A(n571), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U648 ( .A(n572), .B(G143), .Z(G45) );
  XOR2_X1 U649 ( .A(G119), .B(n573), .Z(G21) );
  XNOR2_X1 U650 ( .A(n574), .B(G110), .ZN(G12) );
  INV_X1 U651 ( .A(G475), .ZN(n575) );
  XOR2_X1 U652 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n576) );
  XOR2_X1 U653 ( .A(n577), .B(n576), .Z(n578) );
  XNOR2_X1 U654 ( .A(n579), .B(n578), .ZN(n580) );
  INV_X1 U655 ( .A(n674), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n580), .A2(n588), .ZN(n582) );
  INV_X1 U657 ( .A(KEYINPUT60), .ZN(n581) );
  XNOR2_X1 U658 ( .A(n582), .B(n581), .ZN(G60) );
  NAND2_X1 U659 ( .A1(n592), .A2(G210), .ZN(n587) );
  XNOR2_X1 U660 ( .A(KEYINPUT83), .B(KEYINPUT54), .ZN(n583) );
  XOR2_X1 U661 ( .A(n583), .B(KEYINPUT55), .Z(n584) );
  XNOR2_X1 U662 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U663 ( .A(n587), .B(n586), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n591) );
  XOR2_X1 U665 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n590) );
  XNOR2_X1 U666 ( .A(n591), .B(n590), .ZN(G51) );
  NAND2_X1 U667 ( .A1(n662), .A2(G217), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n593), .B(KEYINPUT123), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n595), .B(n594), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n596), .A2(n674), .ZN(G66) );
  XNOR2_X1 U671 ( .A(G101), .B(n597), .ZN(G3) );
  NOR2_X1 U672 ( .A1(n600), .A2(n610), .ZN(n598) );
  XOR2_X1 U673 ( .A(KEYINPUT114), .B(n598), .Z(n599) );
  XNOR2_X1 U674 ( .A(G104), .B(n599), .ZN(G6) );
  NOR2_X1 U675 ( .A1(n600), .A2(n613), .ZN(n602) );
  XNOR2_X1 U676 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U678 ( .A(G107), .B(n603), .ZN(G9) );
  NOR2_X1 U679 ( .A1(n607), .A2(n613), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n605), .B(n604), .ZN(n606) );
  XOR2_X1 U682 ( .A(G128), .B(n606), .Z(G30) );
  NOR2_X1 U683 ( .A1(n607), .A2(n610), .ZN(n608) );
  XOR2_X1 U684 ( .A(KEYINPUT116), .B(n608), .Z(n609) );
  XNOR2_X1 U685 ( .A(G146), .B(n609), .ZN(G48) );
  NOR2_X1 U686 ( .A1(n612), .A2(n610), .ZN(n611) );
  XOR2_X1 U687 ( .A(G113), .B(n611), .Z(G15) );
  XNOR2_X1 U688 ( .A(G116), .B(KEYINPUT117), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n615), .B(n614), .ZN(G18) );
  XOR2_X1 U691 ( .A(G125), .B(KEYINPUT37), .Z(n616) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(G27) );
  XOR2_X1 U693 ( .A(G134), .B(n618), .Z(G36) );
  INV_X1 U694 ( .A(KEYINPUT81), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n630), .A2(n648), .ZN(n657) );
  INV_X1 U696 ( .A(n620), .ZN(n654) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n628) );
  NOR2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U701 ( .A(KEYINPUT120), .B(n629), .Z(n631) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n651) );
  INV_X1 U703 ( .A(n632), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT49), .B(n635), .Z(n636) );
  NOR2_X1 U706 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT118), .B(n638), .Z(n644) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n641), .B(KEYINPUT50), .ZN(n642) );
  XNOR2_X1 U710 ( .A(KEYINPUT119), .B(n642), .ZN(n643) );
  NOR2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT51), .B(n647), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U715 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U716 ( .A(KEYINPUT52), .B(n652), .Z(n653) );
  NOR2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U718 ( .A1(n655), .A2(G952), .ZN(n656) );
  NAND2_X1 U719 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U720 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U721 ( .A1(n696), .A2(n660), .ZN(n661) );
  XOR2_X1 U722 ( .A(KEYINPUT53), .B(n661), .Z(G75) );
  NAND2_X1 U723 ( .A1(n662), .A2(G469), .ZN(n666) );
  XOR2_X1 U724 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n663) );
  XNOR2_X1 U725 ( .A(n664), .B(n663), .ZN(n665) );
  NOR2_X1 U726 ( .A1(n674), .A2(n667), .ZN(G54) );
  NOR2_X1 U727 ( .A1(n669), .A2(n668), .ZN(n672) );
  XNOR2_X1 U728 ( .A(n670), .B(KEYINPUT122), .ZN(n671) );
  XNOR2_X1 U729 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U730 ( .A1(n674), .A2(n673), .ZN(G63) );
  AND2_X1 U731 ( .A1(n675), .A2(n696), .ZN(n681) );
  NAND2_X1 U732 ( .A1(G953), .A2(G224), .ZN(n676) );
  XNOR2_X1 U733 ( .A(n676), .B(KEYINPUT61), .ZN(n678) );
  NAND2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U735 ( .A(KEYINPUT124), .B(n679), .Z(n680) );
  NOR2_X1 U736 ( .A1(n681), .A2(n680), .ZN(n687) );
  XOR2_X1 U737 ( .A(G101), .B(n682), .Z(n683) );
  XNOR2_X1 U738 ( .A(KEYINPUT125), .B(n683), .ZN(n684) );
  NOR2_X1 U739 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U740 ( .A(n687), .B(n686), .Z(G69) );
  XOR2_X1 U741 ( .A(n689), .B(n688), .Z(n690) );
  XNOR2_X1 U742 ( .A(n691), .B(n690), .ZN(n694) );
  XOR2_X1 U743 ( .A(n694), .B(n693), .Z(n699) );
  XNOR2_X1 U744 ( .A(n695), .B(n699), .ZN(n697) );
  NAND2_X1 U745 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U746 ( .A(KEYINPUT126), .B(n698), .ZN(n704) );
  XOR2_X1 U747 ( .A(G227), .B(n699), .Z(n700) );
  NAND2_X1 U748 ( .A1(n700), .A2(G900), .ZN(n701) );
  NAND2_X1 U749 ( .A1(n701), .A2(G953), .ZN(n702) );
  XOR2_X1 U750 ( .A(KEYINPUT127), .B(n702), .Z(n703) );
  NAND2_X1 U751 ( .A1(n704), .A2(n703), .ZN(G72) );
  XNOR2_X1 U752 ( .A(G140), .B(n705), .ZN(G42) );
  XOR2_X1 U753 ( .A(n706), .B(G122), .Z(G24) );
  XOR2_X1 U754 ( .A(G137), .B(n707), .Z(G39) );
  XOR2_X1 U755 ( .A(n708), .B(G131), .Z(G33) );
endmodule

