

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G651), .A2(n654), .ZN(n657) );
  XOR2_X1 U553 ( .A(KEYINPUT17), .B(n553), .Z(n516) );
  NAND2_X4 U554 ( .A1(n796), .A2(n697), .ZN(n741) );
  XOR2_X1 U555 ( .A(n553), .B(KEYINPUT17), .Z(n900) );
  XNOR2_X1 U556 ( .A(n701), .B(KEYINPUT94), .ZN(n709) );
  OR2_X1 U557 ( .A1(n741), .A2(n698), .ZN(n700) );
  INV_X1 U558 ( .A(n709), .ZN(n710) );
  XNOR2_X1 U559 ( .A(n740), .B(n739), .ZN(n745) );
  NOR2_X1 U560 ( .A1(n825), .A2(n824), .ZN(n827) );
  XNOR2_X1 U561 ( .A(n794), .B(n793), .ZN(n825) );
  XNOR2_X1 U562 ( .A(n522), .B(n521), .ZN(n524) );
  NAND2_X1 U563 ( .A1(n516), .A2(G138), .ZN(n522) );
  XNOR2_X2 U564 ( .A(n526), .B(KEYINPUT64), .ZN(n557) );
  AND2_X1 U565 ( .A1(n556), .A2(n555), .ZN(n517) );
  AND2_X1 U566 ( .A1(n559), .A2(n558), .ZN(n518) );
  NOR2_X1 U567 ( .A1(n773), .A2(n781), .ZN(n519) );
  NAND2_X1 U568 ( .A1(G303), .A2(n744), .ZN(n520) );
  INV_X1 U569 ( .A(KEYINPUT26), .ZN(n702) );
  INV_X1 U570 ( .A(KEYINPUT27), .ZN(n714) );
  XNOR2_X1 U571 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U572 ( .A1(n717), .A2(n716), .ZN(n720) );
  NOR2_X1 U573 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U574 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U575 ( .A(KEYINPUT95), .ZN(n739) );
  NOR2_X1 U576 ( .A1(n761), .A2(n760), .ZN(n763) );
  INV_X1 U577 ( .A(KEYINPUT100), .ZN(n793) );
  NOR2_X2 U578 ( .A1(G2105), .A2(G2104), .ZN(n553) );
  INV_X1 U579 ( .A(KEYINPUT101), .ZN(n826) );
  INV_X1 U580 ( .A(KEYINPUT89), .ZN(n521) );
  OR2_X1 U581 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U582 ( .A(n551), .B(KEYINPUT74), .ZN(n552) );
  XNOR2_X1 U583 ( .A(n540), .B(KEYINPUT68), .ZN(G299) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U585 ( .A1(n897), .A2(G114), .ZN(n523) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n530) );
  INV_X1 U587 ( .A(G2105), .ZN(n525) );
  AND2_X1 U588 ( .A1(n525), .A2(G2104), .ZN(n901) );
  NAND2_X1 U589 ( .A1(G102), .A2(n901), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n525), .A2(G2104), .ZN(n526) );
  NAND2_X1 U591 ( .A1(G126), .A2(n557), .ZN(n527) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(G164) );
  XOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .Z(n654) );
  INV_X1 U595 ( .A(G651), .ZN(n533) );
  NOR2_X2 U596 ( .A1(n654), .A2(n533), .ZN(n666) );
  NAND2_X1 U597 ( .A1(G78), .A2(n666), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G53), .A2(n657), .ZN(n532) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n662) );
  NAND2_X1 U600 ( .A1(G91), .A2(n662), .ZN(n531) );
  NAND2_X1 U601 ( .A1(n532), .A2(n531), .ZN(n537) );
  NOR2_X1 U602 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X2 U603 ( .A(KEYINPUT1), .B(n534), .Z(n659) );
  NAND2_X1 U604 ( .A1(G65), .A2(n659), .ZN(n535) );
  XNOR2_X1 U605 ( .A(KEYINPUT67), .B(n535), .ZN(n536) );
  NOR2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U608 ( .A1(n662), .A2(G89), .ZN(n541) );
  XNOR2_X1 U609 ( .A(KEYINPUT4), .B(n541), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n666), .A2(G76), .ZN(n542) );
  XOR2_X1 U611 ( .A(KEYINPUT73), .B(n542), .Z(n543) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U613 ( .A(n545), .B(KEYINPUT5), .Z(n550) );
  NAND2_X1 U614 ( .A1(G51), .A2(n657), .ZN(n547) );
  NAND2_X1 U615 ( .A1(G63), .A2(n659), .ZN(n546) );
  NAND2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(n552), .ZN(G168) );
  XOR2_X1 U619 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U620 ( .A1(n900), .A2(G137), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G101), .A2(n901), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT23), .B(n554), .Z(n555) );
  NAND2_X1 U623 ( .A1(G113), .A2(n897), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G125), .A2(n557), .ZN(n558) );
  AND2_X1 U625 ( .A1(n517), .A2(n518), .ZN(G160) );
  XOR2_X1 U626 ( .A(G2443), .B(G2451), .Z(n561) );
  XNOR2_X1 U627 ( .A(G2454), .B(G2427), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(n562), .B(G2430), .Z(n564) );
  XNOR2_X1 U630 ( .A(G1341), .B(G1348), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT109), .B(G2435), .Z(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT108), .B(G2438), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U635 ( .A(n568), .B(n567), .Z(n570) );
  XNOR2_X1 U636 ( .A(G2446), .B(KEYINPUT107), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  AND2_X1 U638 ( .A1(n571), .A2(G14), .ZN(G401) );
  NAND2_X1 U639 ( .A1(G52), .A2(n657), .ZN(n573) );
  NAND2_X1 U640 ( .A1(G64), .A2(n659), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G90), .A2(n662), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G77), .A2(n666), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U646 ( .A1(n578), .A2(n577), .ZN(G171) );
  AND2_X1 U647 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U648 ( .A(G82), .ZN(G220) );
  INV_X1 U649 ( .A(G57), .ZN(G237) );
  INV_X1 U650 ( .A(G120), .ZN(G236) );
  INV_X1 U651 ( .A(G108), .ZN(G238) );
  NAND2_X1 U652 ( .A1(G50), .A2(n657), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G75), .A2(n666), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G62), .A2(n659), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT82), .ZN(n584) );
  NAND2_X1 U657 ( .A1(G88), .A2(n662), .ZN(n582) );
  XOR2_X1 U658 ( .A(KEYINPUT83), .B(n582), .Z(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(G166) );
  INV_X1 U661 ( .A(G166), .ZN(G303) );
  NAND2_X1 U662 ( .A1(G7), .A2(G661), .ZN(n587) );
  XNOR2_X1 U663 ( .A(n587), .B(KEYINPUT10), .ZN(n588) );
  XNOR2_X1 U664 ( .A(KEYINPUT70), .B(n588), .ZN(G223) );
  INV_X1 U665 ( .A(G223), .ZN(n850) );
  NAND2_X1 U666 ( .A1(n850), .A2(G567), .ZN(n589) );
  XOR2_X1 U667 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  NAND2_X1 U668 ( .A1(G56), .A2(n659), .ZN(n590) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT14), .ZN(n591) );
  XNOR2_X1 U670 ( .A(KEYINPUT71), .B(n591), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n662), .A2(G81), .ZN(n592) );
  XOR2_X1 U672 ( .A(KEYINPUT12), .B(n592), .Z(n595) );
  NAND2_X1 U673 ( .A1(n666), .A2(G68), .ZN(n593) );
  XOR2_X1 U674 ( .A(KEYINPUT72), .B(n593), .Z(n594) );
  NOR2_X1 U675 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U676 ( .A(KEYINPUT13), .B(n596), .ZN(n597) );
  NOR2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n657), .A2(G43), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n989) );
  INV_X1 U680 ( .A(G860), .ZN(n634) );
  OR2_X1 U681 ( .A1(n989), .A2(n634), .ZN(G153) );
  INV_X1 U682 ( .A(G171), .ZN(G301) );
  NAND2_X1 U683 ( .A1(G868), .A2(G301), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G66), .A2(n659), .ZN(n602) );
  NAND2_X1 U685 ( .A1(G79), .A2(n666), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U687 ( .A1(G54), .A2(n657), .ZN(n604) );
  NAND2_X1 U688 ( .A1(G92), .A2(n662), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U691 ( .A(KEYINPUT15), .B(n607), .Z(n981) );
  INV_X1 U692 ( .A(n981), .ZN(n616) );
  INV_X1 U693 ( .A(G868), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U696 ( .A1(G868), .A2(G286), .ZN(n611) );
  NAND2_X1 U697 ( .A1(G299), .A2(n615), .ZN(n610) );
  NAND2_X1 U698 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U699 ( .A1(G559), .A2(n634), .ZN(n612) );
  XOR2_X1 U700 ( .A(KEYINPUT75), .B(n612), .Z(n613) );
  NAND2_X1 U701 ( .A1(n613), .A2(n981), .ZN(n614) );
  XNOR2_X1 U702 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U704 ( .A(KEYINPUT76), .B(n617), .Z(n618) );
  NOR2_X1 U705 ( .A1(G559), .A2(n618), .ZN(n620) );
  NOR2_X1 U706 ( .A1(G868), .A2(n989), .ZN(n619) );
  NOR2_X1 U707 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G135), .A2(n900), .ZN(n621) );
  XNOR2_X1 U709 ( .A(n621), .B(KEYINPUT78), .ZN(n624) );
  NAND2_X1 U710 ( .A1(G111), .A2(n897), .ZN(n622) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n622), .Z(n623) );
  NAND2_X1 U712 ( .A1(n624), .A2(n623), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n557), .A2(G123), .ZN(n625) );
  XOR2_X1 U714 ( .A(KEYINPUT77), .B(n625), .Z(n626) );
  XNOR2_X1 U715 ( .A(n626), .B(KEYINPUT18), .ZN(n628) );
  NAND2_X1 U716 ( .A1(G99), .A2(n901), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U718 ( .A1(n630), .A2(n629), .ZN(n1010) );
  XNOR2_X1 U719 ( .A(n1010), .B(G2096), .ZN(n632) );
  INV_X1 U720 ( .A(G2100), .ZN(n631) );
  NAND2_X1 U721 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U722 ( .A1(G559), .A2(n981), .ZN(n633) );
  XOR2_X1 U723 ( .A(n989), .B(n633), .Z(n676) );
  NAND2_X1 U724 ( .A1(n634), .A2(n676), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G55), .A2(n657), .ZN(n636) );
  NAND2_X1 U726 ( .A1(G67), .A2(n659), .ZN(n635) );
  NAND2_X1 U727 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U728 ( .A1(G93), .A2(n662), .ZN(n638) );
  NAND2_X1 U729 ( .A1(G80), .A2(n666), .ZN(n637) );
  NAND2_X1 U730 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U731 ( .A1(n640), .A2(n639), .ZN(n678) );
  XOR2_X1 U732 ( .A(n641), .B(n678), .Z(G145) );
  NAND2_X1 U733 ( .A1(G73), .A2(n666), .ZN(n642) );
  XOR2_X1 U734 ( .A(KEYINPUT2), .B(n642), .Z(n645) );
  NAND2_X1 U735 ( .A1(n659), .A2(G61), .ZN(n643) );
  XOR2_X1 U736 ( .A(KEYINPUT80), .B(n643), .Z(n644) );
  NOR2_X1 U737 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U738 ( .A1(n662), .A2(G86), .ZN(n646) );
  NAND2_X1 U739 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U740 ( .A(n648), .B(KEYINPUT81), .ZN(n650) );
  NAND2_X1 U741 ( .A1(G48), .A2(n657), .ZN(n649) );
  NAND2_X1 U742 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U743 ( .A1(G49), .A2(n657), .ZN(n652) );
  NAND2_X1 U744 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U745 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U746 ( .A1(n659), .A2(n653), .ZN(n656) );
  NAND2_X1 U747 ( .A1(n654), .A2(G87), .ZN(n655) );
  NAND2_X1 U748 ( .A1(n656), .A2(n655), .ZN(G288) );
  NAND2_X1 U749 ( .A1(G47), .A2(n657), .ZN(n658) );
  XNOR2_X1 U750 ( .A(n658), .B(KEYINPUT66), .ZN(n661) );
  NAND2_X1 U751 ( .A1(n659), .A2(G60), .ZN(n660) );
  NAND2_X1 U752 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U753 ( .A1(G85), .A2(n662), .ZN(n663) );
  XNOR2_X1 U754 ( .A(KEYINPUT65), .B(n663), .ZN(n664) );
  NOR2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n666), .A2(G72), .ZN(n667) );
  NAND2_X1 U757 ( .A1(n668), .A2(n667), .ZN(G290) );
  XNOR2_X1 U758 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n670) );
  XNOR2_X1 U759 ( .A(G288), .B(KEYINPUT19), .ZN(n669) );
  XNOR2_X1 U760 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U761 ( .A(n678), .B(n671), .ZN(n673) );
  XNOR2_X1 U762 ( .A(G290), .B(G166), .ZN(n672) );
  XNOR2_X1 U763 ( .A(n673), .B(n672), .ZN(n674) );
  XOR2_X1 U764 ( .A(G299), .B(n674), .Z(n675) );
  XNOR2_X1 U765 ( .A(G305), .B(n675), .ZN(n858) );
  XNOR2_X1 U766 ( .A(n676), .B(n858), .ZN(n677) );
  NAND2_X1 U767 ( .A1(n677), .A2(G868), .ZN(n680) );
  OR2_X1 U768 ( .A1(G868), .A2(n678), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U770 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U771 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U772 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U773 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U776 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U777 ( .A1(G238), .A2(G236), .ZN(n685) );
  NAND2_X1 U778 ( .A1(G69), .A2(n685), .ZN(n686) );
  NOR2_X1 U779 ( .A1(n686), .A2(G237), .ZN(n687) );
  XNOR2_X1 U780 ( .A(n687), .B(KEYINPUT87), .ZN(n854) );
  NAND2_X1 U781 ( .A1(n854), .A2(G567), .ZN(n693) );
  NOR2_X1 U782 ( .A1(G220), .A2(G219), .ZN(n688) );
  XOR2_X1 U783 ( .A(KEYINPUT86), .B(n688), .Z(n689) );
  XNOR2_X1 U784 ( .A(n689), .B(KEYINPUT22), .ZN(n690) );
  NOR2_X1 U785 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U786 ( .A1(G96), .A2(n691), .ZN(n855) );
  NAND2_X1 U787 ( .A1(n855), .A2(G2106), .ZN(n692) );
  NAND2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n929) );
  NAND2_X1 U789 ( .A1(G661), .A2(G483), .ZN(n694) );
  XNOR2_X1 U790 ( .A(KEYINPUT88), .B(n694), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n929), .A2(n695), .ZN(n853) );
  NAND2_X1 U792 ( .A1(n853), .A2(G36), .ZN(G176) );
  NOR2_X1 U793 ( .A1(G164), .A2(G1384), .ZN(n796) );
  AND2_X1 U794 ( .A1(G40), .A2(n518), .ZN(n696) );
  NAND2_X1 U795 ( .A1(n696), .A2(n517), .ZN(n795) );
  INV_X1 U796 ( .A(n795), .ZN(n697) );
  INV_X1 U797 ( .A(G2067), .ZN(n698) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n741), .ZN(n699) );
  NAND2_X1 U799 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U800 ( .A1(n616), .A2(n709), .ZN(n708) );
  INV_X1 U801 ( .A(n741), .ZN(n713) );
  AND2_X1 U802 ( .A1(n713), .A2(G1996), .ZN(n703) );
  XNOR2_X1 U803 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U804 ( .A1(n741), .A2(G1341), .ZN(n704) );
  NAND2_X1 U805 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U806 ( .A1(n989), .A2(n706), .ZN(n707) );
  NAND2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n710), .A2(n981), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n713), .A2(G2072), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G1956), .A2(n741), .ZN(n716) );
  NOR2_X1 U812 ( .A1(G299), .A2(n720), .ZN(n718) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U814 ( .A1(G299), .A2(n720), .ZN(n721) );
  XOR2_X1 U815 ( .A(KEYINPUT28), .B(n721), .Z(n722) );
  XNOR2_X1 U816 ( .A(n724), .B(KEYINPUT29), .ZN(n729) );
  INV_X1 U817 ( .A(n741), .ZN(n725) );
  OR2_X1 U818 ( .A1(n725), .A2(G1961), .ZN(n727) );
  XNOR2_X1 U819 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NAND2_X1 U820 ( .A1(n725), .A2(n957), .ZN(n726) );
  NAND2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n733) );
  NAND2_X1 U822 ( .A1(G171), .A2(n733), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n738) );
  NAND2_X1 U824 ( .A1(G8), .A2(n741), .ZN(n773) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n773), .ZN(n752) );
  NOR2_X1 U826 ( .A1(G2084), .A2(n741), .ZN(n748) );
  NOR2_X1 U827 ( .A1(n752), .A2(n748), .ZN(n730) );
  NAND2_X1 U828 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  NOR2_X1 U830 ( .A1(G168), .A2(n732), .ZN(n735) );
  NOR2_X1 U831 ( .A1(G171), .A2(n733), .ZN(n734) );
  XOR2_X1 U832 ( .A(KEYINPUT31), .B(n736), .Z(n737) );
  NAND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n749) );
  NAND2_X1 U834 ( .A1(n749), .A2(G286), .ZN(n740) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n773), .ZN(n743) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n741), .ZN(n742) );
  NOR2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n745), .A2(n520), .ZN(n746) );
  NAND2_X1 U839 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U840 ( .A(KEYINPUT32), .B(n747), .ZN(n776) );
  NAND2_X1 U841 ( .A1(G8), .A2(n748), .ZN(n754) );
  BUF_X1 U842 ( .A(n749), .Z(n750) );
  INV_X1 U843 ( .A(n750), .ZN(n751) );
  NOR2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n774) );
  AND2_X1 U846 ( .A1(n774), .A2(n773), .ZN(n755) );
  AND2_X1 U847 ( .A1(n776), .A2(n755), .ZN(n761) );
  INV_X1 U848 ( .A(n773), .ZN(n759) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n756) );
  XNOR2_X1 U850 ( .A(n756), .B(KEYINPUT98), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n757), .A2(G8), .ZN(n758) );
  NOR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  INV_X1 U853 ( .A(KEYINPUT99), .ZN(n762) );
  XNOR2_X1 U854 ( .A(n763), .B(n762), .ZN(n767) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U856 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  OR2_X1 U857 ( .A1(n773), .A2(n765), .ZN(n766) );
  AND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n792) );
  INV_X1 U859 ( .A(KEYINPUT33), .ZN(n771) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n779) );
  INV_X1 U861 ( .A(n779), .ZN(n768) );
  NOR2_X1 U862 ( .A1(KEYINPUT96), .A2(n768), .ZN(n769) );
  NOR2_X1 U863 ( .A1(n773), .A2(n769), .ZN(n770) );
  NOR2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n788) );
  NAND2_X1 U865 ( .A1(n779), .A2(KEYINPUT33), .ZN(n772) );
  NAND2_X1 U866 ( .A1(KEYINPUT96), .A2(n772), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n976) );
  AND2_X1 U868 ( .A1(n519), .A2(n976), .ZN(n777) );
  AND2_X1 U869 ( .A1(n774), .A2(n777), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n786) );
  INV_X1 U871 ( .A(n777), .ZN(n780) );
  NOR2_X1 U872 ( .A1(G1971), .A2(G303), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n977) );
  NOR2_X1 U874 ( .A1(n780), .A2(n977), .ZN(n784) );
  INV_X1 U875 ( .A(n781), .ZN(n782) );
  AND2_X1 U876 ( .A1(n782), .A2(KEYINPUT33), .ZN(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n790) );
  XOR2_X1 U880 ( .A(KEYINPUT97), .B(G1981), .Z(n789) );
  XNOR2_X1 U881 ( .A(G305), .B(n789), .ZN(n991) );
  OR2_X1 U882 ( .A1(n790), .A2(n991), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n844) );
  NAND2_X1 U885 ( .A1(G140), .A2(n900), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G104), .A2(n901), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(n799), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G116), .A2(n897), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G128), .A2(n557), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT91), .B(n802), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT35), .B(n803), .ZN(n804) );
  NOR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n806), .ZN(n919) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n831) );
  NOR2_X1 U897 ( .A1(n919), .A2(n831), .ZN(n1023) );
  NAND2_X1 U898 ( .A1(n844), .A2(n1023), .ZN(n841) );
  XOR2_X1 U899 ( .A(n844), .B(KEYINPUT93), .Z(n823) );
  NAND2_X1 U900 ( .A1(G107), .A2(n897), .ZN(n808) );
  NAND2_X1 U901 ( .A1(G119), .A2(n557), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n900), .A2(G131), .ZN(n809) );
  XOR2_X1 U904 ( .A(KEYINPUT92), .B(n809), .Z(n810) );
  NOR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n901), .A2(G95), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n908) );
  NAND2_X1 U908 ( .A1(G1991), .A2(n908), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G141), .A2(n900), .ZN(n815) );
  NAND2_X1 U910 ( .A1(G117), .A2(n897), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n901), .A2(G105), .ZN(n816) );
  XOR2_X1 U913 ( .A(KEYINPUT38), .B(n816), .Z(n817) );
  NOR2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U915 ( .A1(G129), .A2(n557), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n909) );
  NAND2_X1 U917 ( .A1(G1996), .A2(n909), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n1012) );
  NAND2_X1 U919 ( .A1(n823), .A2(n1012), .ZN(n836) );
  NAND2_X1 U920 ( .A1(n841), .A2(n836), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n827), .B(n826), .ZN(n830) );
  XNOR2_X1 U922 ( .A(KEYINPUT90), .B(G1986), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n828), .B(G290), .ZN(n988) );
  NAND2_X1 U924 ( .A1(n988), .A2(n844), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n847) );
  AND2_X1 U926 ( .A1(n831), .A2(n919), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(KEYINPUT105), .ZN(n1020) );
  NOR2_X1 U928 ( .A1(G1986), .A2(G290), .ZN(n834) );
  NOR2_X1 U929 ( .A1(n908), .A2(G1991), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n833), .B(KEYINPUT102), .ZN(n1011) );
  NOR2_X1 U931 ( .A1(n834), .A2(n1011), .ZN(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT103), .B(n835), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(n838) );
  OR2_X1 U934 ( .A1(n909), .A2(G1996), .ZN(n1015) );
  NAND2_X1 U935 ( .A1(n838), .A2(n1015), .ZN(n840) );
  XOR2_X1 U936 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n1020), .A2(n843), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U941 ( .A1(n847), .A2(n846), .ZN(n849) );
  XNOR2_X1 U942 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n848) );
  XNOR2_X1 U943 ( .A(n849), .B(n848), .ZN(G329) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U946 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(G188) );
  XOR2_X1 U949 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U953 ( .A(G286), .B(KEYINPUT117), .ZN(n857) );
  XNOR2_X1 U954 ( .A(G171), .B(n981), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n860) );
  XOR2_X1 U956 ( .A(n989), .B(n858), .Z(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(n861) );
  NOR2_X1 U958 ( .A1(G37), .A2(n861), .ZN(G397) );
  XOR2_X1 U959 ( .A(G2100), .B(G2096), .Z(n863) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(G2678), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U962 ( .A(KEYINPUT43), .B(G2090), .Z(n865) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2072), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U966 ( .A(G2078), .B(G2084), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(G227) );
  XOR2_X1 U968 ( .A(G1956), .B(G1961), .Z(n871) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1991), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U971 ( .A(G1966), .B(G1971), .Z(n873) );
  XNOR2_X1 U972 ( .A(G1981), .B(G1976), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U975 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(G2474), .B(n878), .ZN(n879) );
  XOR2_X1 U978 ( .A(n879), .B(G1996), .Z(G229) );
  NAND2_X1 U979 ( .A1(n557), .A2(G124), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n880), .B(KEYINPUT44), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G112), .A2(n897), .ZN(n881) );
  XOR2_X1 U982 ( .A(KEYINPUT113), .B(n881), .Z(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n900), .A2(G136), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(KEYINPUT112), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G100), .A2(n901), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(G162) );
  NAND2_X1 U989 ( .A1(G139), .A2(n900), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G103), .A2(n901), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U992 ( .A(KEYINPUT114), .B(n891), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G115), .A2(n897), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G127), .A2(n557), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n1003) );
  NAND2_X1 U998 ( .A1(G118), .A2(n897), .ZN(n899) );
  NAND2_X1 U999 ( .A1(G130), .A2(n557), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n900), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n901), .ZN(n902) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT45), .B(n904), .Z(n905) );
  NOR2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n1003), .B(n907), .ZN(n918) );
  XNOR2_X1 U1007 ( .A(n1010), .B(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1009 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G162), .B(KEYINPUT48), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1012 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1013 ( .A(G164), .B(G160), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1016 ( .A(n920), .B(n919), .Z(n921) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT116), .B(n922), .ZN(G395) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n929), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n924), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(n927), .A2(G395), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(n928), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1026 ( .A(G308), .ZN(G225) );
  INV_X1 U1027 ( .A(n929), .ZN(G319) );
  INV_X1 U1028 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1029 ( .A(KEYINPUT125), .B(G1966), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(n930), .B(G21), .ZN(n948) );
  XOR2_X1 U1031 ( .A(G1348), .B(KEYINPUT59), .Z(n931) );
  XNOR2_X1 U1032 ( .A(G4), .B(n931), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G20), .B(G1956), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(KEYINPUT60), .ZN(n946) );
  XOR2_X1 U1040 ( .A(G1986), .B(G24), .Z(n942) );
  XNOR2_X1 U1041 ( .A(G1976), .B(G23), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n939) );
  NOR2_X1 U1043 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(n943), .B(KEYINPUT126), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(KEYINPUT58), .B(n944), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(G5), .B(G1961), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(KEYINPUT61), .B(n951), .ZN(n953) );
  INV_X1 U1052 ( .A(G16), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n974) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n954) );
  NOR2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n963) );
  XOR2_X1 U1057 ( .A(G1991), .B(G25), .Z(n956) );
  NAND2_X1 U1058 ( .A1(n956), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(n957), .B(G27), .ZN(n959) );
  XOR2_X1 U1060 ( .A(G1996), .B(G32), .Z(n958) );
  NAND2_X1 U1061 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1062 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1064 ( .A(n964), .B(KEYINPUT53), .ZN(n967) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(KEYINPUT122), .B(G2090), .ZN(n968) );
  XNOR2_X1 U1069 ( .A(G35), .B(n968), .ZN(n969) );
  NOR2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n1033) );
  INV_X1 U1071 ( .A(n1033), .ZN(n972) );
  NOR2_X1 U1072 ( .A1(G29), .A2(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n1002) );
  XOR2_X1 U1075 ( .A(G16), .B(KEYINPUT56), .Z(n1000) );
  XNOR2_X1 U1076 ( .A(G171), .B(G1961), .ZN(n986) );
  INV_X1 U1077 ( .A(G1971), .ZN(n975) );
  NOR2_X1 U1078 ( .A1(G166), .A2(n975), .ZN(n979) );
  NAND2_X1 U1079 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1080 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1081 ( .A(KEYINPUT124), .B(n980), .Z(n984) );
  XNOR2_X1 U1082 ( .A(G1348), .B(n981), .ZN(n982) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n982), .ZN(n983) );
  NOR2_X1 U1084 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1085 ( .A1(n986), .A2(n985), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1956), .B(G299), .ZN(n987) );
  NOR2_X1 U1087 ( .A1(n988), .A2(n987), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n989), .B(G1341), .ZN(n994) );
  XOR2_X1 U1089 ( .A(G1966), .B(G168), .Z(n990) );
  NOR2_X1 U1090 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1091 ( .A(KEYINPUT57), .B(n992), .ZN(n993) );
  NOR2_X1 U1092 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1093 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1094 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1032) );
  XNOR2_X1 U1097 ( .A(G2072), .B(n1003), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(n1004), .B(KEYINPUT121), .ZN(n1006) );
  XOR2_X1 U1099 ( .A(G2078), .B(G164), .Z(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1101 ( .A(KEYINPUT50), .B(n1007), .Z(n1026) );
  XNOR2_X1 U1102 ( .A(G160), .B(G2084), .ZN(n1008) );
  XNOR2_X1 U1103 ( .A(n1008), .B(KEYINPUT119), .ZN(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G162), .B(G2090), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1109 ( .A(KEYINPUT51), .B(n1017), .Z(n1018) );
  NOR2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(KEYINPUT120), .B(n1024), .Z(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  INV_X1 U1116 ( .A(KEYINPUT55), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1036) );
  NAND2_X1 U1120 ( .A1(KEYINPUT55), .A2(n1033), .ZN(n1034) );
  NAND2_X1 U1121 ( .A1(G11), .A2(n1034), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1123 ( .A(n1037), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

