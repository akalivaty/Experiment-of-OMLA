//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT67), .Z(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  AOI211_X1 g0026(.A(new_n213), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n243), .A2(G1), .A3(G13), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G226), .A3(new_n250), .ZN(new_n251));
  OR2_X1    g0051(.A1(new_n251), .A2(KEYINPUT73), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(KEYINPUT73), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n249), .A2(G232), .A3(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n244), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n244), .A3(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n244), .A2(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(G238), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT13), .B1(new_n259), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT13), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n257), .B1(new_n252), .B2(new_n253), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n267), .C1(new_n271), .C2(new_n244), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(KEYINPUT74), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n259), .A2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT74), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n270), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(G169), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT14), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(KEYINPUT76), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n273), .A2(new_n276), .A3(G169), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n269), .A2(G179), .A3(new_n272), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT77), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT77), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n269), .A2(new_n272), .A3(new_n285), .A4(G179), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n222), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G50), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n292), .A2(new_n293), .B1(new_n223), .B2(G68), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n223), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT11), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n290), .B1(new_n260), .B2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n303), .A2(KEYINPUT12), .A3(G68), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT12), .B1(new_n303), .B2(G68), .ZN(new_n305));
  AOI22_X1  g0105(.A1(G68), .A2(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n288), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n273), .A2(G200), .A3(new_n276), .ZN(new_n310));
  INV_X1    g0110(.A(new_n307), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n269), .A2(G190), .A3(new_n272), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n303), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n293), .ZN(new_n317));
  INV_X1    g0117(.A(new_n302), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n293), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n291), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT8), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n320), .B1(new_n295), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n319), .B1(new_n327), .B2(new_n290), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT9), .Z(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G222), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n249), .A2(G1698), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n334), .B1(new_n296), .B2(new_n249), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n244), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n264), .B1(G226), .B2(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G190), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n329), .B(new_n343), .C1(new_n344), .C2(new_n342), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT72), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT10), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n345), .B(new_n347), .Z(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n328), .B1(new_n341), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n321), .A2(new_n292), .B1(new_n223), .B2(new_n296), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT15), .B(G87), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n356), .A2(new_n357), .B1(new_n359), .B2(new_n295), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n356), .A2(new_n357), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n290), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT71), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n303), .A2(G77), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n302), .B2(G77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n266), .A2(G244), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n249), .A2(G232), .A3(new_n250), .ZN(new_n369));
  INV_X1    g0169(.A(G107), .ZN(new_n370));
  INV_X1    g0170(.A(G238), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n369), .B1(new_n370), .B2(new_n249), .C1(new_n336), .C2(new_n371), .ZN(new_n372));
  AOI211_X1 g0172(.A(new_n264), .B(new_n368), .C1(new_n372), .C2(new_n338), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n367), .B(new_n374), .C1(new_n344), .C2(new_n373), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(G169), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n352), .B2(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n366), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n335), .A2(G1698), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n330), .B2(new_n331), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  OAI211_X1 g0183(.A(G226), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT78), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n380), .B(new_n385), .C1(new_n331), .C2(new_n330), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n338), .ZN(new_n388));
  INV_X1    g0188(.A(G232), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n263), .B1(new_n389), .B2(new_n265), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n352), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n387), .B2(new_n338), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(G169), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n290), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n332), .B2(new_n223), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n248), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G68), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n324), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n202), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n291), .A2(G159), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n395), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n247), .A2(new_n223), .A3(new_n248), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n400), .B1(new_n410), .B2(new_n397), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n402), .A2(new_n403), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n326), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n318), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n326), .A2(new_n303), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n406), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT18), .B1(new_n394), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n416), .ZN(new_n419));
  INV_X1    g0219(.A(new_n412), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT16), .B1(new_n399), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n290), .B1(new_n411), .B2(new_n404), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n388), .A2(new_n391), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n349), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n423), .A2(new_n425), .A3(new_n426), .A4(new_n392), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(G200), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n393), .A2(G190), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n417), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n417), .A2(new_n429), .A3(KEYINPUT17), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n379), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n315), .A2(new_n348), .A3(new_n355), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  AND2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G257), .A3(new_n244), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(G274), .A3(new_n244), .A4(new_n440), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G244), .B(new_n250), .C1(new_n330), .C2(new_n331), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n250), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AOI211_X1 g0254(.A(KEYINPUT81), .B(new_n447), .C1(new_n454), .C2(new_n338), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n338), .ZN(new_n457));
  INV_X1    g0257(.A(new_n447), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G190), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n292), .A2(new_n296), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n370), .A2(KEYINPUT6), .A3(G97), .ZN(new_n464));
  XNOR2_X1  g0264(.A(G97), .B(G107), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT6), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(new_n223), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n370), .B1(new_n410), .B2(new_n397), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n290), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n396), .B2(new_n398), .ZN(new_n472));
  AND2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n370), .A2(KEYINPUT6), .A3(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n462), .B1(new_n477), .B2(G20), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n290), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n260), .A2(G33), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n395), .A2(KEYINPUT80), .A3(new_n303), .A4(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n303), .A2(new_n483), .A3(new_n222), .A4(new_n289), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G97), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(G97), .B2(new_n316), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n457), .A2(new_n458), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G200), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n461), .A2(new_n482), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n457), .A2(new_n352), .A3(new_n458), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n482), .B2(new_n490), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n349), .B1(new_n455), .B2(new_n459), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G190), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n244), .A2(G274), .A3(new_n440), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n260), .A2(G45), .ZN(new_n504));
  AND2_X1   g0304(.A1(G33), .A2(G41), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n504), .B(G250), .C1(new_n505), .C2(new_n222), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G238), .B(new_n250), .C1(new_n330), .C2(new_n331), .ZN(new_n508));
  OAI211_X1 g0308(.A(G244), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n502), .B(new_n507), .C1(new_n338), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n338), .ZN(new_n513));
  INV_X1    g0313(.A(new_n507), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n344), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n358), .A2(new_n303), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n223), .B1(new_n256), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n474), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n223), .B(G68), .C1(new_n330), .C2(new_n331), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n518), .B1(new_n295), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n517), .B1(new_n526), .B2(new_n290), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n484), .A2(new_n487), .A3(G87), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n507), .B1(new_n511), .B2(new_n338), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n484), .A2(new_n487), .A3(new_n358), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n352), .A2(new_n530), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n513), .A2(new_n514), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n349), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n516), .A2(new_n529), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n493), .A2(new_n498), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(KEYINPUT82), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n453), .B(new_n223), .C1(G33), .C2(new_n524), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n539), .B(new_n290), .C1(new_n223), .C2(G116), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT20), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n316), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n485), .B2(new_n542), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n443), .A2(new_n244), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G270), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n547), .A2(new_n446), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n249), .A2(G264), .A3(G1698), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n249), .A2(G257), .A3(new_n250), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n332), .A2(G303), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n552), .A2(new_n553), .A3(new_n338), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n552), .B2(new_n338), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n545), .B1(G200), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n502), .B2(new_n556), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT84), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n548), .B(G179), .C1(new_n554), .C2(new_n555), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n541), .A2(new_n544), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n547), .A2(new_n446), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n552), .A2(new_n338), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT83), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n552), .A2(new_n553), .A3(new_n338), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(new_n545), .A3(KEYINPUT84), .A4(G179), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G169), .B1(new_n541), .B2(new_n544), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT21), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n556), .A2(new_n545), .A3(new_n572), .A4(G169), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n558), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n546), .A2(G264), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n249), .A2(G257), .A3(G1698), .ZN(new_n577));
  INV_X1    g0377(.A(G294), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n246), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT86), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n333), .A2(new_n580), .A3(G250), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n249), .A2(G250), .A3(new_n250), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT86), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n446), .B(new_n576), .C1(new_n584), .C2(new_n244), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n349), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n581), .A2(new_n583), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n338), .B1(new_n587), .B2(new_n579), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(new_n352), .A3(new_n446), .A4(new_n576), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n249), .A2(new_n223), .A3(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT22), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n249), .A2(new_n593), .A3(new_n223), .A4(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n370), .A3(G20), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT85), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n596), .B2(new_n370), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n597), .A2(new_n598), .B1(new_n601), .B2(G20), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n590), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n595), .A2(new_n590), .A3(new_n603), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n395), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n484), .A2(new_n487), .A3(G107), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n303), .A2(G107), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT25), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n586), .B(new_n589), .C1(new_n607), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n585), .A2(G200), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n588), .A2(G190), .A3(new_n446), .A4(new_n576), .ZN(new_n614));
  INV_X1    g0414(.A(new_n606), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n290), .B1(new_n615), .B2(new_n604), .ZN(new_n616));
  INV_X1    g0416(.A(new_n611), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n613), .A2(new_n614), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT87), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT87), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n612), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n575), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n438), .A2(new_n501), .A3(new_n538), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n355), .ZN(new_n625));
  INV_X1    g0425(.A(new_n378), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n309), .B1(new_n313), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n418), .A2(KEYINPUT91), .A3(new_n427), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT91), .B1(new_n418), .B2(new_n427), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n627), .A2(new_n435), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n630), .B2(new_n348), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n533), .A2(KEYINPUT88), .A3(new_n349), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT88), .B1(new_n533), .B2(new_n349), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n532), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n480), .B1(new_n479), .B2(new_n290), .ZN(new_n635));
  AOI211_X1 g0435(.A(KEYINPUT79), .B(new_n395), .C1(new_n472), .C2(new_n478), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n490), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n497), .A2(new_n494), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .A3(new_n535), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT90), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n516), .A2(new_n529), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n498), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n612), .B(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n569), .A2(new_n574), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n634), .A2(new_n643), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n618), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n653), .A2(new_n498), .A3(new_n493), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n631), .B1(new_n437), .B2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n260), .A2(new_n223), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI211_X1 g0464(.A(new_n561), .B(new_n664), .C1(new_n569), .C2(new_n574), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT92), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(KEYINPUT92), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n575), .B1(new_n545), .B2(new_n663), .ZN(new_n668));
  OAI211_X1 g0468(.A(G330), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n620), .A2(new_n622), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n663), .B1(new_n607), .B2(new_n611), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n612), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n663), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n649), .A2(new_n663), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n650), .A2(new_n663), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n670), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n211), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n474), .A2(new_n520), .A3(new_n542), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n685), .A2(new_n260), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n226), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT28), .Z(new_n689));
  AOI21_X1  g0489(.A(new_n663), .B1(new_n647), .B2(new_n655), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT95), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n642), .B1(new_n638), .B2(new_n652), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n496), .A2(new_n642), .A3(new_n497), .A4(new_n535), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n634), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n498), .B2(new_n644), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(KEYINPUT95), .A3(new_n634), .A4(new_n695), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n612), .A2(new_n569), .A3(new_n574), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n653), .A2(new_n700), .A3(new_n498), .A4(new_n493), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n691), .B1(new_n702), .B2(new_n664), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n692), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  XOR2_X1   g0505(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n706));
  NOR3_X1   g0506(.A1(new_n567), .A2(G179), .A3(new_n530), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT94), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n585), .A2(new_n708), .A3(new_n491), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n585), .B2(new_n491), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n560), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n530), .B(new_n576), .C1(new_n584), .C2(new_n244), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n460), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n460), .A2(new_n712), .A3(new_n714), .A4(KEYINPUT30), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n711), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n663), .ZN(new_n720));
  MUX2_X1   g0520(.A(new_n706), .B(KEYINPUT31), .S(new_n720), .Z(new_n721));
  NAND4_X1  g0521(.A1(new_n623), .A2(new_n501), .A3(new_n538), .A4(new_n664), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n705), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n704), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n689), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT98), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(G1), .B(G13), .C1(new_n223), .C2(G169), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT99), .Z(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n684), .A2(new_n249), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n241), .A2(new_n439), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n738), .B(new_n739), .C1(new_n439), .C2(new_n226), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n211), .A2(G355), .A3(new_n249), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G116), .B2(new_n211), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n736), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n209), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n260), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n685), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT96), .Z(new_n748));
  NOR3_X1   g0548(.A1(new_n502), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n223), .ZN(new_n750));
  NAND2_X1  g0550(.A1(G20), .A2(G179), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(new_n344), .A3(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n524), .B1(new_n753), .B2(new_n400), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT100), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n223), .A2(G179), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT32), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n756), .A2(new_n502), .A3(G200), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n760), .B(new_n249), .C1(new_n370), .C2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n751), .A2(new_n502), .A3(new_n344), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n751), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n757), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n293), .B1(new_n766), .B2(new_n296), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n751), .A2(new_n502), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n502), .A2(new_n344), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n756), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n769), .A2(new_n324), .B1(new_n771), .B2(new_n520), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n758), .A2(KEYINPUT32), .A3(new_n759), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n762), .A2(new_n767), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n758), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n775), .A2(G329), .B1(new_n768), .B2(G322), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n249), .B1(new_n763), .B2(G326), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n750), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G294), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n753), .A2(new_n781), .B1(new_n761), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n771), .A2(new_n784), .B1(new_n766), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n755), .A2(new_n774), .B1(new_n780), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n743), .B(new_n748), .C1(new_n788), .C2(new_n734), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n732), .ZN(new_n791));
  INV_X1    g0591(.A(new_n669), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n747), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n790), .A2(new_n705), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  OAI21_X1  g0596(.A(new_n375), .B1(new_n367), .B2(new_n664), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n378), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n626), .A2(new_n664), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n690), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT102), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n690), .A2(new_n801), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n723), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT103), .ZN(new_n810));
  INV_X1    g0610(.A(new_n747), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n724), .B1(new_n806), .B2(new_n807), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT103), .B1(new_n813), .B2(new_n747), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(new_n723), .C2(new_n808), .ZN(new_n815));
  INV_X1    g0615(.A(new_n748), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G137), .A2(new_n763), .B1(new_n752), .B2(G150), .ZN(new_n817));
  INV_X1    g0617(.A(G143), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n818), .B2(new_n769), .C1(new_n759), .C2(new_n766), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n249), .B1(new_n771), .B2(new_n293), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n761), .A2(new_n400), .B1(new_n758), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(G58), .C2(new_n779), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n332), .B1(new_n771), .B2(new_n370), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT101), .ZN(new_n829));
  INV_X1    g0629(.A(new_n761), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(G87), .B1(new_n768), .B2(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n753), .A2(new_n782), .B1(new_n766), .B2(new_n542), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G97), .B2(new_n779), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n775), .A2(G311), .B1(G303), .B2(new_n763), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n829), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n734), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n735), .A2(new_n728), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n816), .B(new_n836), .C1(new_n296), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n801), .B2(new_n729), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n815), .A2(new_n839), .ZN(G384));
  OR2_X1    g0640(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(G116), .A4(new_n224), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  OAI211_X1 g0644(.A(new_n226), .B(G77), .C1(new_n324), .C2(new_n400), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n201), .A2(G68), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n260), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n849));
  INV_X1    g0649(.A(new_n706), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n719), .B2(new_n663), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n722), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n438), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT108), .ZN(new_n855));
  INV_X1    g0655(.A(new_n661), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n423), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n431), .B(new_n857), .C1(new_n417), .C2(new_n394), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(new_n857), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n435), .B2(new_n428), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n858), .B(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n433), .A2(new_n434), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n628), .B2(new_n629), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n860), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n865), .B1(new_n868), .B2(KEYINPUT106), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT106), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT107), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT91), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n428), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n418), .A2(KEYINPUT91), .A3(new_n427), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n435), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT106), .B1(new_n878), .B2(new_n857), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n871), .A3(new_n859), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n307), .A2(new_n663), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n308), .A2(new_n886), .A3(new_n313), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n307), .B(new_n663), .C1(new_n288), .C2(new_n314), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND4_X1   g0689(.A1(KEYINPUT40), .A2(new_n889), .A3(new_n853), .A4(new_n801), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n859), .B2(new_n861), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n863), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT105), .A3(new_n862), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n800), .B1(new_n852), .B2(new_n722), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n889), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n884), .A2(new_n890), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n855), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n855), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(G330), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n802), .A2(new_n799), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n896), .A3(new_n889), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n876), .A2(new_n877), .A3(new_n661), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n880), .A2(new_n873), .A3(new_n881), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n862), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n910), .B2(new_n882), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n863), .A2(new_n908), .A3(new_n892), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n308), .A2(new_n663), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n906), .B(new_n907), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n438), .B1(new_n692), .B2(new_n703), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n631), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n904), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n260), .B2(new_n744), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n904), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n848), .B1(new_n922), .B2(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n637), .A2(new_n663), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n499), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n638), .A2(new_n663), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n679), .A3(new_n681), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT45), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n928), .B1(new_n679), .B2(new_n681), .ZN(new_n933));
  NOR2_X1   g0733(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n682), .A2(new_n928), .A3(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n678), .A2(KEYINPUT111), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n931), .B1(new_n936), .B2(new_n937), .C1(KEYINPUT111), .C2(new_n678), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n681), .B1(new_n675), .B2(new_n680), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n669), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n704), .A3(new_n724), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT112), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n725), .A2(new_n944), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT112), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(new_n949), .A3(new_n940), .A4(new_n941), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n725), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n685), .B(new_n952), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n745), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n928), .A2(new_n670), .A3(new_n680), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n493), .A2(new_n673), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n663), .B1(new_n957), .B2(new_n498), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n955), .B2(KEYINPUT42), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n529), .A2(new_n664), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n652), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n634), .A2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n956), .A2(new_n959), .B1(KEYINPUT43), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n677), .A2(new_n928), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n954), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n736), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n738), .A2(new_n234), .B1(new_n211), .B2(new_n359), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n748), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n771), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT113), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n830), .A2(G97), .B1(new_n768), .B2(G303), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n979), .B(new_n332), .C1(new_n980), .C2(new_n758), .ZN(new_n981));
  INV_X1    g0781(.A(new_n766), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n982), .A2(G283), .B1(G294), .B2(new_n752), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n785), .B2(new_n764), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n974), .A2(new_n975), .B1(new_n370), .B2(new_n750), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n775), .A2(G137), .B1(G143), .B2(new_n763), .ZN(new_n987));
  INV_X1    g0787(.A(new_n201), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n982), .A2(new_n988), .B1(G150), .B2(new_n768), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n249), .B1(new_n753), .B2(new_n759), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n750), .A2(new_n400), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n761), .A2(new_n296), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n771), .A2(new_n324), .ZN(new_n994));
  NOR4_X1   g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n978), .A2(new_n986), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n734), .B1(new_n996), .B2(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n972), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n961), .A2(new_n732), .A3(new_n962), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n969), .A2(new_n1001), .ZN(G387));
  NAND2_X1  g0802(.A1(new_n725), .A2(new_n944), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n946), .A3(new_n685), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n779), .A2(G283), .B1(new_n973), .B2(G294), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G322), .A2(new_n763), .B1(new_n752), .B2(G311), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n784), .B2(new_n766), .C1(new_n980), .C2(new_n769), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT115), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT49), .Z(new_n1013));
  AOI21_X1  g0813(.A(new_n249), .B1(new_n775), .B2(G326), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n542), .B2(new_n761), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT116), .Z(new_n1016));
  NOR2_X1   g0816(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n771), .A2(new_n296), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G159), .B2(new_n763), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n332), .B1(new_n830), .B2(G97), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G150), .A2(new_n775), .B1(new_n982), .B2(G68), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n359), .A2(new_n750), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G50), .B2(new_n768), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT114), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1025), .C1(new_n414), .C2(new_n752), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n735), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n970), .B1(G107), .B2(new_n684), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n231), .A2(new_n439), .A3(new_n249), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n321), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT50), .B1(new_n321), .B2(G50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n686), .B1(new_n1033), .B2(new_n332), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n211), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n816), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n676), .B2(new_n732), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n945), .B2(new_n746), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1004), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT117), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT117), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1004), .A2(new_n1042), .A3(new_n1039), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(G393));
  AOI22_X1  g0844(.A1(G317), .A2(new_n763), .B1(new_n768), .B2(G311), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT52), .Z(new_n1046));
  AOI22_X1  g0846(.A1(G283), .A2(new_n973), .B1(new_n775), .B2(G322), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n982), .A2(G294), .B1(G303), .B2(new_n752), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n332), .B1(new_n761), .B2(new_n370), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G116), .B2(new_n779), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G150), .A2(new_n763), .B1(new_n768), .B2(G159), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT51), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n750), .A2(new_n296), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n332), .B(new_n1054), .C1(G87), .C2(new_n830), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n753), .A2(new_n201), .B1(new_n758), .B2(new_n818), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n771), .A2(new_n400), .B1(new_n766), .B2(new_n321), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n734), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n738), .A2(new_n238), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G97), .B2(new_n684), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n816), .B(new_n1060), .C1(new_n736), .C2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n928), .B2(new_n731), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n938), .B(new_n677), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n745), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n947), .A2(new_n950), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n685), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(new_n946), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(G390));
  AOI22_X1  g0871(.A1(new_n690), .A2(new_n798), .B1(new_n626), .B2(new_n664), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n889), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n916), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT39), .B1(new_n874), .B2(new_n883), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n912), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n723), .A2(new_n801), .A3(new_n889), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT118), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n915), .B1(new_n874), .B2(new_n883), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n702), .A2(new_n664), .A3(new_n798), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n799), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n889), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1078), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n916), .C1(new_n910), .C2(new_n882), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1084), .A2(KEYINPUT118), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1076), .B(new_n1077), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1079), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(KEYINPUT118), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1087), .A2(new_n1088), .B1(new_n914), .B2(new_n1074), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n897), .A2(new_n889), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1090), .A2(new_n705), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n705), .B1(new_n852), .B2(new_n722), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n438), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n631), .A2(new_n918), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n889), .B1(new_n723), .B2(new_n801), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n905), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n801), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1073), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1077), .A2(new_n1100), .A3(new_n799), .A4(new_n1080), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1096), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1086), .B(new_n1102), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n685), .A3(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1093), .A2(new_n745), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n816), .B1(new_n326), .B2(new_n837), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n973), .A2(G150), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G159), .B2(new_n779), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n982), .A2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n775), .A2(G125), .B1(new_n752), .B2(G137), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n764), .A2(new_n1116), .B1(new_n769), .B2(new_n824), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n332), .B(new_n1117), .C1(new_n988), .C2(new_n830), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .A4(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n332), .B1(new_n771), .B2(new_n520), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT119), .Z(new_n1121));
  AOI22_X1  g0921(.A1(new_n982), .A2(G97), .B1(G107), .B2(new_n752), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n775), .A2(G294), .B1(new_n768), .B2(G116), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n764), .A2(new_n782), .B1(new_n761), .B2(new_n400), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n1054), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1075), .A2(new_n912), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1108), .B1(new_n734), .B2(new_n1127), .C1(new_n1128), .C2(new_n729), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1106), .A2(new_n1107), .A3(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(new_n1096), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1105), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n348), .A2(new_n355), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n328), .A2(new_n661), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n348), .B(new_n355), .C1(new_n328), .C2(new_n661), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n900), .B2(G330), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n890), .B1(new_n882), .B2(new_n910), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n898), .A2(new_n899), .ZN(new_n1146));
  AND4_X1   g0946(.A1(G330), .A2(new_n1145), .A3(new_n1146), .A4(new_n1143), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n917), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n906), .A2(new_n907), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n915), .B2(new_n1128), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n900), .A2(G330), .A3(new_n1143), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1145), .A2(new_n1146), .A3(G330), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1143), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1133), .B1(new_n1148), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT121), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1132), .A2(new_n1156), .A3(KEYINPUT121), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1105), .A2(new_n1131), .B1(new_n1155), .B2(new_n1148), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n685), .B1(new_n1162), .B2(KEYINPUT57), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1143), .A2(new_n729), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n1116), .A2(new_n769), .B1(new_n753), .B2(new_n824), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n982), .A2(G137), .B1(new_n763), .B2(G125), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n771), .B2(new_n1112), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G150), .C2(new_n779), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT59), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  INV_X1    g0973(.A(G41), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n246), .B(new_n1174), .C1(new_n761), .C2(new_n759), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G124), .B2(new_n775), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n753), .A2(new_n524), .B1(new_n761), .B2(new_n324), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n332), .A2(new_n1174), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1178), .A2(new_n992), .A3(new_n1018), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n768), .A2(G107), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT120), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n763), .A2(G116), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G283), .A2(new_n775), .B1(new_n982), .B2(new_n358), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1179), .B(new_n293), .C1(G33), .C2(G41), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1177), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n735), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n811), .B(new_n1191), .C1(new_n201), .C2(new_n837), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1165), .A2(new_n746), .B1(new_n1166), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1164), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G375));
  AND2_X1   g0996(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1096), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n953), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1103), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1073), .A2(new_n728), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n982), .A2(G107), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n768), .A2(G283), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n542), .B2(new_n753), .C1(new_n784), .C2(new_n758), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n973), .A2(G97), .B1(new_n763), .B2(G294), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1209), .A2(new_n1023), .A3(new_n993), .A4(new_n249), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n982), .A2(G150), .B1(G137), .B2(new_n768), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1113), .A2(new_n752), .B1(G132), .B2(new_n763), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G159), .A2(new_n973), .B1(new_n775), .B2(G128), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n332), .B1(new_n830), .B2(G58), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n293), .C2(new_n750), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1207), .A2(new_n1210), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(new_n734), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n816), .B(new_n1219), .C1(new_n400), .C2(new_n837), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1201), .A2(new_n746), .B1(new_n1202), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1200), .A2(new_n1221), .ZN(G381));
  INV_X1    g1022(.A(new_n1001), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n954), .B2(new_n968), .ZN(new_n1224));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1041), .A2(new_n795), .A3(new_n1043), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1195), .A2(new_n1224), .A3(new_n1225), .A4(new_n1227), .ZN(G407));
  INV_X1    g1028(.A(G213), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(G343), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1195), .A2(new_n1225), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(G213), .A3(new_n1231), .ZN(G409));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n815), .A2(new_n1233), .A3(new_n839), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n815), .B2(new_n839), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1197), .A2(KEYINPUT60), .A3(new_n1096), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n685), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1103), .A2(KEYINPUT60), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1198), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1221), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1234), .A2(new_n1235), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1198), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n685), .A3(new_n1236), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1221), .C1(KEYINPUT122), .C2(G384), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1193), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1162), .A2(new_n1199), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1225), .B1(new_n1194), .B2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1230), .B(new_n1245), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT123), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT63), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1230), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(KEYINPUT123), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT125), .B1(new_n1224), .B2(G390), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1043), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1042), .B1(new_n1004), .B2(new_n1039), .ZN(new_n1259));
  OAI21_X1  g1059(.A(G396), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1226), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT124), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1226), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1224), .A2(G390), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1223), .B(new_n1070), .C1(new_n954), .C2(new_n968), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1257), .A2(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(new_n1070), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1260), .A2(new_n1226), .A3(new_n1263), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1263), .B1(new_n1260), .B2(new_n1226), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1224), .A2(G390), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1272), .A3(KEYINPUT125), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1268), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1252), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1230), .A2(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1241), .A2(new_n1244), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1276), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1251), .A2(new_n1256), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1252), .A2(new_n1286), .A3(new_n1253), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1252), .B2(new_n1282), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1287), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1268), .A2(new_n1274), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1285), .B1(new_n1291), .B2(new_n1293), .ZN(G405));
  AND2_X1   g1094(.A1(new_n1253), .A2(KEYINPUT127), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1292), .B(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1246), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1195), .A2(G378), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1298), .A2(new_n1297), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(G402));
endmodule


