//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n462), .B2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n488), .A2(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(G62), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n497), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n504), .A2(G651), .B1(G50), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n500), .B(new_n502), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT69), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(G88), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(new_n512), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n513), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n520), .B(new_n522), .C1(new_n528), .C2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n519), .A2(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n503), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(G52), .B2(new_n507), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n519), .A2(G81), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n503), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(G43), .B2(new_n507), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  XOR2_X1   g123(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n549));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n524), .A2(new_n553), .B1(KEYINPUT73), .B2(KEYINPUT9), .ZN(new_n554));
  NOR2_X1   g129(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n507), .B(G53), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(KEYINPUT74), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G651), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n512), .A2(new_n516), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n562), .A2(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n508), .A2(new_n517), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(G303));
  NAND2_X1  g148(.A1(new_n519), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n507), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n500), .A2(new_n502), .A3(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n507), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n512), .A2(G86), .A3(new_n516), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n507), .A2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n564), .B2(new_n585), .C1(new_n566), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n519), .A2(new_n589), .A3(G92), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n503), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT10), .B1(new_n566), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT76), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n588), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n588), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n568), .B1(new_n561), .B2(new_n560), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n598), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n477), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  NAND2_X1  g188(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n613), .B(new_n614), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n475), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n477), .A2(G135), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  OAI211_X1 g196(.A(new_n615), .B(new_n621), .C1(KEYINPUT77), .C2(G2100), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT78), .Z(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2438), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n633), .B(new_n634), .Z(new_n635));
  AND2_X1   g210(.A1(new_n635), .A2(G14), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT79), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT18), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n638), .B(KEYINPUT80), .Z(new_n646));
  INV_X1    g221(.A(new_n642), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n638), .B(KEYINPUT17), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n644), .B1(new_n645), .B2(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT81), .B(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  AND2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT82), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT83), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n670), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  OAI21_X1  g249(.A(KEYINPUT92), .B1(G5), .B2(G16), .ZN(new_n675));
  OR3_X1    g250(.A1(KEYINPUT92), .A2(G5), .A3(G16), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n675), .B(new_n676), .C1(G301), .C2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G1961), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(KEYINPUT23), .A3(G20), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n682));
  INV_X1    g257(.A(G20), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G16), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n684), .C1(new_n602), .C2(new_n677), .ZN(new_n685));
  INV_X1    g260(.A(G1956), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G35), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G162), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT29), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n687), .A2(new_n688), .B1(G2090), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n680), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n677), .A2(G19), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n545), .B2(new_n677), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1341), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G11), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(G28), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(G28), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(new_n702), .A3(new_n689), .ZN(new_n703));
  OAI221_X1 g278(.A(new_n703), .B1(new_n689), .B2(new_n620), .C1(new_n692), .C2(G2090), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n689), .A2(G26), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT87), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  OR2_X1    g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT86), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n475), .A2(G128), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n477), .A2(G140), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2067), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n689), .A2(G27), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G164), .B2(new_n689), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(G2078), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n704), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n695), .A2(new_n698), .A3(new_n699), .A4(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n687), .A2(new_n688), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n692), .A2(G2090), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT93), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n477), .A2(G139), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT88), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  AOI22_X1  g302(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT89), .Z(new_n729));
  OAI211_X1 g304(.A(new_n725), .B(new_n727), .C1(new_n462), .C2(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G33), .B(new_n730), .S(G29), .Z(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G2072), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n679), .B2(new_n678), .ZN(new_n733));
  NAND2_X1  g308(.A1(G168), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G21), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(KEYINPUT91), .A3(new_n736), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n740), .A2(new_n741), .B1(new_n731), .B2(G2072), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n723), .A2(new_n733), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n689), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n689), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2084), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n720), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G32), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n486), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n753), .A2(new_n462), .B1(new_n475), .B2(G129), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT90), .Z(new_n759));
  AOI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(G16), .A2(G23), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G288), .B2(new_n677), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT33), .B(G1976), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n677), .A2(G22), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G166), .B2(new_n677), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n677), .A2(G6), .ZN(new_n772));
  INV_X1    g347(.A(G305), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n677), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT32), .B(G1981), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n766), .A2(new_n770), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n689), .A2(G25), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n475), .A2(G119), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT84), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n477), .A2(G131), .ZN(new_n781));
  NOR2_X1   g356(.A1(G95), .A2(G2105), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n689), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT35), .B(G1991), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G24), .B(G290), .S(G16), .Z(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1986), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n777), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT85), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n777), .A2(new_n788), .A3(new_n793), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n766), .A2(new_n770), .A3(new_n776), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n796), .B1(new_n795), .B2(new_n798), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n750), .B(new_n762), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n677), .A2(G4), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n598), .B2(new_n677), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1348), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n717), .A2(G2078), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n802), .A2(new_n805), .A3(new_n807), .ZN(G311));
  NOR2_X1   g383(.A1(new_n720), .A2(new_n749), .ZN(new_n809));
  INV_X1    g384(.A(new_n743), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n801), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n799), .ZN(new_n813));
  INV_X1    g388(.A(new_n805), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n813), .A2(new_n814), .A3(new_n806), .A4(new_n762), .ZN(G150));
  XNOR2_X1  g390(.A(KEYINPUT95), .B(G93), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n519), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n507), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n564), .ZN(new_n821));
  OAI21_X1  g396(.A(G860), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n598), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT39), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n826));
  INV_X1    g401(.A(new_n821), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n817), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n817), .A2(new_n827), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n545), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n817), .A2(new_n827), .A3(new_n826), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n832), .A2(new_n828), .A3(new_n544), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n825), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n823), .B1(new_n838), .B2(G860), .ZN(G145));
  XOR2_X1   g414(.A(new_n785), .B(new_n612), .Z(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n489), .A2(new_n841), .A3(new_n493), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n489), .B2(new_n493), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n485), .B(new_n487), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n620), .B(G160), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n481), .ZN(new_n848));
  AOI22_X1  g423(.A1(G130), .A2(new_n475), .B1(new_n477), .B2(G142), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT98), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT98), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n851), .B(new_n852), .C1(G118), .C2(new_n462), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n713), .B(new_n854), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n848), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n758), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n730), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n759), .B2(new_n730), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n846), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n856), .A2(new_n859), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n845), .A3(new_n860), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g443(.A(G288), .B(G290), .Z(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g447(.A1(G166), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n571), .A2(KEYINPUT100), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n773), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(G305), .A3(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(G288), .B(G290), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n871), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n876), .A2(new_n879), .A3(KEYINPUT101), .A4(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n607), .B(new_n834), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n597), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n602), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n888), .A2(KEYINPUT99), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT99), .B1(new_n888), .B2(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n887), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n887), .A2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n818), .A2(new_n821), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(G868), .B2(new_n904), .ZN(G295));
  OAI21_X1  g480(.A(new_n903), .B1(G868), .B2(new_n904), .ZN(G331));
  NAND2_X1  g481(.A1(G171), .A2(G286), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n526), .B(new_n527), .ZN(new_n908));
  NAND4_X1  g483(.A1(G301), .A2(new_n908), .A3(new_n520), .A4(new_n522), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n831), .B2(new_n833), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n829), .A2(new_n545), .A3(new_n830), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n544), .B1(new_n832), .B2(new_n828), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n907), .A4(new_n909), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n892), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n895), .A2(new_n911), .A3(new_n896), .A4(new_n914), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(KEYINPUT104), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n911), .A2(new_n914), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n897), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n881), .A2(new_n882), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n916), .B1(new_n918), .B2(new_n892), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n883), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n864), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT105), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n922), .A2(new_n927), .A3(new_n864), .A4(new_n924), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(KEYINPUT43), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n921), .B1(new_n917), .B2(new_n920), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(G37), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n922), .A2(new_n933), .A3(new_n864), .A4(new_n924), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n932), .B2(new_n933), .ZN(new_n937));
  XOR2_X1   g512(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n941));
  INV_X1    g516(.A(G1981), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n581), .A2(new_n582), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n581), .B2(new_n582), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G8), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n494), .A2(KEYINPUT97), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n489), .A2(new_n841), .A3(new_n493), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n488), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n467), .A2(new_n468), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G2105), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n472), .A2(new_n462), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n955), .A2(new_n956), .A3(G40), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n948), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n943), .ZN(new_n959));
  INV_X1    g534(.A(new_n944), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(KEYINPUT49), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(KEYINPUT110), .B(new_n941), .C1(new_n943), .C2(new_n944), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n947), .A2(new_n958), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n574), .A2(G1976), .A3(new_n575), .A4(new_n576), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT52), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(G288), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n958), .A3(new_n964), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n963), .A2(new_n966), .A3(KEYINPUT114), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(G303), .B2(G8), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n571), .A2(new_n572), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT75), .B1(new_n508), .B2(new_n517), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n975), .B(G8), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT106), .B(G1384), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n844), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n488), .B2(new_n494), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n957), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n769), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n955), .A2(new_n956), .A3(G40), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n993));
  NAND3_X1  g568(.A1(new_n844), .A2(new_n985), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(G2090), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n990), .B(new_n998), .C1(G2090), .C2(new_n995), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n981), .A2(new_n997), .A3(G8), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n993), .B1(new_n844), .B2(new_n985), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n991), .ZN(new_n1003));
  INV_X1    g578(.A(G2090), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT113), .B(new_n957), .C1(new_n953), .C2(new_n993), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n990), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT55), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n979), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT45), .B(new_n985), .C1(new_n488), .C2(new_n494), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n957), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n488), .B1(new_n949), .B2(new_n950), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n987), .B1(new_n1017), .B2(G1384), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1966), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n992), .A2(new_n994), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G286), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n974), .A2(new_n1000), .A3(new_n1013), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n972), .A2(new_n973), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(KEYINPUT115), .A3(new_n1000), .A4(new_n1023), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n997), .A2(G8), .A3(new_n999), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n970), .B1(new_n1031), .B2(new_n1012), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT63), .A3(new_n1000), .A4(new_n1023), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1003), .A2(new_n1006), .A3(new_n1005), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n686), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n558), .B(new_n565), .C1(new_n567), .C2(new_n566), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n1037), .B2(KEYINPUT116), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n562), .A2(new_n569), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(KEYINPUT57), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT56), .B(G2072), .Z(new_n1042));
  OR2_X1    g617(.A1(new_n989), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1036), .B2(new_n1043), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1348), .B1(new_n992), .B2(new_n994), .ZN(new_n1046));
  NOR4_X1   g621(.A1(new_n1017), .A2(new_n991), .A3(G1384), .A4(G2067), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n597), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT61), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1036), .A2(new_n1041), .A3(new_n1051), .A4(new_n1043), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(KEYINPUT119), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1046), .A2(new_n1055), .A3(new_n1047), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n890), .B1(new_n1056), .B2(KEYINPUT120), .ZN(new_n1057));
  INV_X1    g632(.A(G1348), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n995), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1047), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(KEYINPUT60), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n597), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1057), .A2(new_n1063), .B1(KEYINPUT120), .B2(new_n1056), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1048), .A2(KEYINPUT60), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1052), .B(new_n1054), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  OR3_X1    g642(.A1(new_n989), .A2(new_n1067), .A3(G1996), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n985), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(new_n991), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1067), .B1(new_n989), .B2(G1996), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n544), .B1(new_n1074), .B2(KEYINPUT59), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(KEYINPUT118), .A3(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1073), .B(new_n1075), .C1(new_n1074), .C2(KEYINPUT59), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1050), .B1(new_n1066), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1028), .A2(new_n1000), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n989), .B2(G2078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n995), .A2(new_n679), .ZN(new_n1086));
  INV_X1    g661(.A(G2078), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1016), .A2(new_n1018), .A3(KEYINPUT53), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n1089), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT124), .B1(new_n1089), .B2(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1017), .A2(new_n982), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n957), .B1(new_n1095), .B2(KEYINPUT45), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n984), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n844), .A2(new_n983), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n991), .B1(new_n1099), .B2(new_n987), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT53), .B(new_n1087), .C1(new_n1100), .C2(KEYINPUT122), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1087), .A2(KEYINPUT53), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1100), .A2(KEYINPUT122), .B1(KEYINPUT45), .B2(new_n1095), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT123), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1094), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1102), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(KEYINPUT123), .A3(new_n1106), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1093), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1110), .B1(new_n1113), .B2(G301), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1092), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G286), .A2(G8), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1022), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT51), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT45), .B1(new_n844), .B2(new_n985), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n736), .B1(new_n1123), .B2(new_n1015), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(G2084), .B2(new_n995), .ZN(new_n1125));
  OAI211_X1 g700(.A(G8), .B(new_n1122), .C1(new_n1125), .C2(G286), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(G8), .A3(G286), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1121), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(G301), .B(new_n1094), .C1(new_n1103), .C2(new_n1107), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1089), .A2(G171), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1132), .B2(new_n1083), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1081), .A2(new_n1082), .A3(new_n1115), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1128), .B2(KEYINPUT62), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1121), .A2(new_n1126), .A3(new_n1136), .A4(new_n1127), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1135), .A2(new_n1000), .A3(new_n1028), .A4(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1000), .A2(new_n970), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G288), .A2(G1976), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT112), .Z(new_n1141));
  AND2_X1   g716(.A1(new_n1141), .A2(new_n963), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n943), .B(KEYINPUT111), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n958), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1138), .A2(new_n1139), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1034), .A2(new_n1134), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1099), .A2(new_n987), .A3(new_n957), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(G1996), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n759), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT107), .Z(new_n1150));
  INV_X1    g725(.A(new_n1147), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n713), .B(G2067), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n758), .A2(G1996), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n785), .B(new_n787), .Z(new_n1155));
  OAI211_X1 g730(.A(new_n1150), .B(new_n1154), .C1(new_n1147), .C2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(G1986), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1146), .A2(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1156), .A2(KEYINPUT127), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1147), .A2(G1986), .A3(G290), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT48), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1156), .A2(KEYINPUT127), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1148), .A2(KEYINPUT46), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1151), .B1(new_n1152), .B2(new_n758), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1148), .A2(KEYINPUT46), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT47), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n785), .A2(new_n787), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT126), .Z(new_n1172));
  OAI22_X1  g747(.A1(new_n1170), .A2(new_n1172), .B1(G2067), .B2(new_n713), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1173), .B2(new_n1151), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1164), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1159), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g751(.A(G227), .B1(new_n635), .B2(G14), .ZN(new_n1178));
  AND2_X1   g752(.A1(new_n867), .A2(new_n1178), .ZN(new_n1179));
  AND4_X1   g753(.A1(new_n460), .A2(new_n937), .A3(new_n1179), .A4(new_n673), .ZN(G308));
  NAND4_X1  g754(.A1(new_n937), .A2(new_n1179), .A3(new_n460), .A4(new_n673), .ZN(G225));
endmodule


