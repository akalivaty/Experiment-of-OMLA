

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n752), .B(n751), .ZN(n753) );
  BUF_X1 U550 ( .A(n652), .Z(n516) );
  XNOR2_X1 U551 ( .A(n543), .B(KEYINPUT65), .ZN(n652) );
  AND2_X1 U552 ( .A1(n697), .A2(n696), .ZN(n701) );
  INV_X1 U553 ( .A(n693), .ZN(n723) );
  INV_X1 U554 ( .A(n723), .ZN(n743) );
  NOR2_X1 U555 ( .A1(n754), .A2(n753), .ZN(n803) );
  AND2_X1 U556 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U557 ( .A1(n807), .A2(n806), .ZN(n514) );
  BUF_X1 U558 ( .A(n652), .Z(n515) );
  NOR2_X2 U559 ( .A1(n539), .A2(n538), .ZN(G160) );
  AND2_X2 U560 ( .A1(n527), .A2(G2104), .ZN(n876) );
  XNOR2_X1 U561 ( .A(KEYINPUT0), .B(G543), .ZN(n541) );
  NOR2_X4 U562 ( .A1(G651), .A2(n649), .ZN(n586) );
  INV_X1 U563 ( .A(n975), .ZN(n756) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n720) );
  INV_X1 U565 ( .A(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U566 ( .A1(n757), .A2(n756), .ZN(n758) );
  INV_X1 U567 ( .A(G2104), .ZN(n522) );
  XOR2_X1 U568 ( .A(KEYINPUT31), .B(n735), .Z(n517) );
  OR2_X1 U569 ( .A1(n761), .A2(KEYINPUT33), .ZN(n518) );
  OR2_X1 U570 ( .A1(n795), .A2(n799), .ZN(n519) );
  OR2_X2 U571 ( .A1(n542), .A2(n547), .ZN(n543) );
  AND2_X1 U572 ( .A1(n796), .A2(n519), .ZN(n520) );
  INV_X1 U573 ( .A(KEYINPUT26), .ZN(n694) );
  INV_X1 U574 ( .A(KEYINPUT100), .ZN(n698) );
  INV_X1 U575 ( .A(KEYINPUT101), .ZN(n708) );
  NOR2_X1 U576 ( .A1(n731), .A2(G168), .ZN(n734) );
  NOR2_X1 U577 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U578 ( .A(n721), .B(n720), .ZN(n728) );
  NAND2_X1 U579 ( .A1(G8), .A2(n743), .ZN(n799) );
  INV_X1 U580 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U581 ( .A1(G160), .A2(G40), .ZN(n763) );
  XNOR2_X1 U582 ( .A(n523), .B(KEYINPUT64), .ZN(n524) );
  NOR2_X1 U583 ( .A1(n582), .A2(n581), .ZN(n583) );
  BUF_X1 U584 ( .A(n532), .Z(n610) );
  NOR2_X1 U585 ( .A1(G2104), .A2(n527), .ZN(n879) );
  INV_X1 U586 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n876), .A2(G102), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT17), .B(n524), .ZN(n532) );
  NAND2_X1 U590 ( .A1(G138), .A2(n610), .ZN(n525) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U592 ( .A1(G126), .A2(n879), .ZN(n529) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U594 ( .A1(G114), .A2(n880), .ZN(n528) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U597 ( .A1(G137), .A2(n532), .ZN(n535) );
  NAND2_X1 U598 ( .A1(G101), .A2(n876), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U601 ( .A1(G125), .A2(n879), .ZN(n537) );
  NAND2_X1 U602 ( .A1(G113), .A2(n880), .ZN(n536) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U604 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U605 ( .A1(n654), .A2(G89), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT4), .ZN(n545) );
  INV_X1 U607 ( .A(n541), .ZN(n542) );
  INV_X1 U608 ( .A(G651), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G76), .A2(n516), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT5), .ZN(n553) );
  NOR2_X1 U612 ( .A1(G543), .A2(n547), .ZN(n548) );
  XOR2_X2 U613 ( .A(KEYINPUT1), .B(n548), .Z(n657) );
  NAND2_X1 U614 ( .A1(G63), .A2(n657), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT0), .B(G543), .Z(n649) );
  NAND2_X1 U616 ( .A1(G51), .A2(n586), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U621 ( .A1(G65), .A2(n657), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT70), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G78), .A2(n516), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT69), .B(n556), .Z(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G53), .A2(n586), .ZN(n559) );
  XNOR2_X1 U627 ( .A(KEYINPUT71), .B(n559), .ZN(n560) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n654), .A2(G91), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(G299) );
  NAND2_X1 U631 ( .A1(n516), .A2(G77), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT68), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G90), .A2(n654), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT9), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G64), .A2(n657), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G52), .A2(n586), .ZN(n570) );
  XNOR2_X1 U639 ( .A(KEYINPUT67), .B(n570), .ZN(n571) );
  NOR2_X1 U640 ( .A1(n572), .A2(n571), .ZN(G171) );
  AND2_X1 U641 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U642 ( .A1(n657), .A2(G56), .ZN(n573) );
  XNOR2_X1 U643 ( .A(n573), .B(KEYINPUT14), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G43), .A2(n586), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n515), .A2(G68), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n654), .A2(G81), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U650 ( .A(KEYINPUT74), .B(n579), .Z(n580) );
  XNOR2_X1 U651 ( .A(KEYINPUT13), .B(n580), .ZN(n581) );
  XNOR2_X1 U652 ( .A(KEYINPUT75), .B(n583), .ZN(n691) );
  BUF_X1 U653 ( .A(n691), .Z(n969) );
  INV_X1 U654 ( .A(G860), .ZN(n622) );
  OR2_X1 U655 ( .A1(n969), .A2(n622), .ZN(G153) );
  INV_X1 U656 ( .A(G57), .ZN(G237) );
  XOR2_X1 U657 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U658 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U660 ( .A(G223), .ZN(n829) );
  NAND2_X1 U661 ( .A1(n829), .A2(G567), .ZN(n585) );
  XOR2_X1 U662 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U663 ( .A1(G171), .A2(G868), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G92), .A2(n654), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n586), .A2(G54), .ZN(n587) );
  XOR2_X1 U666 ( .A(KEYINPUT77), .B(n587), .Z(n589) );
  NAND2_X1 U667 ( .A1(n516), .A2(G79), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U669 ( .A(KEYINPUT78), .B(n590), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n657), .A2(G66), .ZN(n591) );
  XOR2_X1 U671 ( .A(KEYINPUT76), .B(n591), .Z(n592) );
  NOR2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U674 ( .A(n596), .B(KEYINPUT15), .Z(n597) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT79), .ZN(n700) );
  BUF_X1 U676 ( .A(n700), .Z(n981) );
  INV_X1 U677 ( .A(G868), .ZN(n671) );
  NAND2_X1 U678 ( .A1(n981), .A2(n671), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U680 ( .A(KEYINPUT80), .B(n600), .Z(G284) );
  NOR2_X1 U681 ( .A1(G286), .A2(n671), .ZN(n602) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U683 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n622), .A2(G559), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n603), .A2(n981), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  INV_X1 U687 ( .A(G559), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n605), .A2(n981), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n606), .A2(G868), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n969), .A2(n671), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U692 ( .A1(n879), .A2(G123), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G135), .A2(n610), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U696 ( .A(n613), .B(KEYINPUT81), .ZN(n615) );
  NAND2_X1 U697 ( .A1(G99), .A2(n876), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n880), .A2(G111), .ZN(n616) );
  XOR2_X1 U700 ( .A(KEYINPUT82), .B(n616), .Z(n617) );
  NOR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n925) );
  XNOR2_X1 U702 ( .A(n925), .B(G2096), .ZN(n620) );
  INV_X1 U703 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(G156) );
  NAND2_X1 U705 ( .A1(G559), .A2(n981), .ZN(n621) );
  XOR2_X1 U706 ( .A(n969), .B(n621), .Z(n668) );
  NAND2_X1 U707 ( .A1(n622), .A2(n668), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G67), .A2(n657), .ZN(n624) );
  NAND2_X1 U709 ( .A1(G55), .A2(n586), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G93), .A2(n654), .ZN(n625) );
  XNOR2_X1 U712 ( .A(KEYINPUT83), .B(n625), .ZN(n626) );
  NOR2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n516), .A2(G80), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n672) );
  XNOR2_X1 U716 ( .A(n630), .B(n672), .ZN(G145) );
  NAND2_X1 U717 ( .A1(G60), .A2(n657), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G47), .A2(n586), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n516), .A2(G72), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n654), .A2(G85), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U724 ( .A(KEYINPUT66), .B(n637), .Z(G290) );
  NAND2_X1 U725 ( .A1(G88), .A2(n654), .ZN(n638) );
  XOR2_X1 U726 ( .A(KEYINPUT86), .B(n638), .Z(n643) );
  NAND2_X1 U727 ( .A1(G62), .A2(n657), .ZN(n640) );
  NAND2_X1 U728 ( .A1(G50), .A2(n586), .ZN(n639) );
  NAND2_X1 U729 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U730 ( .A(KEYINPUT85), .B(n641), .Z(n642) );
  NOR2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n516), .A2(G75), .ZN(n644) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  NAND2_X1 U735 ( .A1(G49), .A2(n586), .ZN(n647) );
  NAND2_X1 U736 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U738 ( .A1(n657), .A2(n648), .ZN(n651) );
  NAND2_X1 U739 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U740 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U741 ( .A1(G73), .A2(n516), .ZN(n653) );
  XNOR2_X1 U742 ( .A(n653), .B(KEYINPUT2), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G48), .A2(n586), .ZN(n656) );
  NAND2_X1 U744 ( .A1(G86), .A2(n654), .ZN(n655) );
  NAND2_X1 U745 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U746 ( .A1(n657), .A2(G61), .ZN(n658) );
  XOR2_X1 U747 ( .A(KEYINPUT84), .B(n658), .Z(n659) );
  NOR2_X1 U748 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n662), .A2(n661), .ZN(G305) );
  XNOR2_X1 U750 ( .A(KEYINPUT19), .B(G288), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n663), .B(n672), .ZN(n664) );
  XNOR2_X1 U752 ( .A(G166), .B(n664), .ZN(n666) );
  INV_X1 U753 ( .A(G299), .ZN(n968) );
  XNOR2_X1 U754 ( .A(G305), .B(n968), .ZN(n665) );
  XNOR2_X1 U755 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U756 ( .A(G290), .B(n667), .ZN(n901) );
  XOR2_X1 U757 ( .A(n668), .B(n901), .Z(n669) );
  XNOR2_X1 U758 ( .A(KEYINPUT87), .B(n669), .ZN(n670) );
  NOR2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n674) );
  NOR2_X1 U760 ( .A1(G868), .A2(n672), .ZN(n673) );
  NOR2_X1 U761 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U768 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  XNOR2_X1 U769 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U770 ( .A1(G219), .A2(G220), .ZN(n679) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U772 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U773 ( .A1(G96), .A2(n681), .ZN(n835) );
  AND2_X1 U774 ( .A1(G2106), .A2(n835), .ZN(n686) );
  NAND2_X1 U775 ( .A1(G69), .A2(G120), .ZN(n682) );
  NOR2_X1 U776 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U777 ( .A1(G108), .A2(n683), .ZN(n834) );
  NAND2_X1 U778 ( .A1(G567), .A2(n834), .ZN(n684) );
  XOR2_X1 U779 ( .A(KEYINPUT88), .B(n684), .Z(n685) );
  NOR2_X1 U780 ( .A1(n686), .A2(n685), .ZN(G319) );
  INV_X1 U781 ( .A(G319), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n833) );
  NAND2_X1 U784 ( .A1(n833), .A2(G36), .ZN(G176) );
  XNOR2_X1 U785 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n828) );
  NOR2_X1 U786 ( .A1(G164), .A2(G1384), .ZN(n764) );
  XOR2_X1 U787 ( .A(KEYINPUT94), .B(n763), .Z(n689) );
  NAND2_X1 U788 ( .A1(n764), .A2(n689), .ZN(n693) );
  NOR2_X1 U789 ( .A1(G1966), .A2(n799), .ZN(n741) );
  AND2_X1 U790 ( .A1(n693), .A2(G1341), .ZN(n690) );
  NOR2_X1 U791 ( .A1(n691), .A2(n690), .ZN(n697) );
  INV_X1 U792 ( .A(G1996), .ZN(n692) );
  NOR2_X1 U793 ( .A1(n693), .A2(n692), .ZN(n695) );
  XNOR2_X1 U794 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X2 U795 ( .A1(n700), .A2(n701), .ZN(n699) );
  XNOR2_X1 U796 ( .A(n699), .B(n698), .ZN(n707) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n723), .A2(G1348), .ZN(n703) );
  NOR2_X1 U799 ( .A1(G2067), .A2(n743), .ZN(n702) );
  NOR2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U803 ( .A(n709), .B(n708), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G2072), .A2(n723), .ZN(n711) );
  XNOR2_X1 U805 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n710) );
  XNOR2_X1 U806 ( .A(n711), .B(n710), .ZN(n713) );
  XNOR2_X1 U807 ( .A(G1956), .B(KEYINPUT99), .ZN(n998) );
  NOR2_X1 U808 ( .A1(n723), .A2(n998), .ZN(n712) );
  NOR2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n716), .A2(n968), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n716), .A2(n968), .ZN(n717) );
  XOR2_X1 U813 ( .A(n717), .B(KEYINPUT28), .Z(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n721) );
  XOR2_X1 U815 ( .A(G2078), .B(KEYINPUT25), .Z(n722) );
  XNOR2_X1 U816 ( .A(KEYINPUT96), .B(n722), .ZN(n952) );
  NAND2_X1 U817 ( .A1(n952), .A2(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G1961), .A2(n743), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U820 ( .A(n726), .B(KEYINPUT97), .ZN(n732) );
  NAND2_X1 U821 ( .A1(G171), .A2(n732), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n736) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n743), .ZN(n738) );
  NOR2_X1 U824 ( .A1(n741), .A2(n738), .ZN(n729) );
  NAND2_X1 U825 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U826 ( .A(n730), .B(KEYINPUT30), .ZN(n731) );
  NOR2_X1 U827 ( .A1(G171), .A2(n732), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n736), .A2(n517), .ZN(n737) );
  XNOR2_X1 U829 ( .A(n737), .B(KEYINPUT102), .ZN(n742) );
  NAND2_X1 U830 ( .A1(G8), .A2(n738), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n742), .A2(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n754) );
  NAND2_X1 U833 ( .A1(n742), .A2(G286), .ZN(n750) );
  INV_X1 U834 ( .A(G8), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n799), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n746), .A2(G303), .ZN(n747) );
  OR2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  AND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n752) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n755), .B(KEYINPUT103), .ZN(n757) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NOR2_X1 U844 ( .A1(n803), .A2(n758), .ZN(n760) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n979) );
  INV_X1 U846 ( .A(n799), .ZN(n805) );
  NAND2_X1 U847 ( .A1(n979), .A2(n805), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U849 ( .A(KEYINPUT104), .B(G1981), .Z(n762) );
  XNOR2_X1 U850 ( .A(G305), .B(n762), .ZN(n989) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n823) );
  NAND2_X1 U852 ( .A1(n879), .A2(G119), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G131), .A2(n610), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G95), .A2(n876), .ZN(n768) );
  NAND2_X1 U856 ( .A1(G107), .A2(n880), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n887) );
  NAND2_X1 U859 ( .A1(G1991), .A2(n887), .ZN(n771) );
  XOR2_X1 U860 ( .A(KEYINPUT91), .B(n771), .Z(n782) );
  NAND2_X1 U861 ( .A1(G105), .A2(n876), .ZN(n772) );
  XOR2_X1 U862 ( .A(KEYINPUT38), .B(n772), .Z(n778) );
  NAND2_X1 U863 ( .A1(n880), .A2(G117), .ZN(n773) );
  XNOR2_X1 U864 ( .A(n773), .B(KEYINPUT92), .ZN(n775) );
  NAND2_X1 U865 ( .A1(G129), .A2(n879), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U867 ( .A(KEYINPUT93), .B(n776), .Z(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U869 ( .A1(G141), .A2(n610), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n891) );
  NAND2_X1 U871 ( .A1(G1996), .A2(n891), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n816) );
  INV_X1 U873 ( .A(n816), .ZN(n794) );
  XNOR2_X1 U874 ( .A(G2067), .B(KEYINPUT37), .ZN(n783) );
  XOR2_X1 U875 ( .A(n783), .B(KEYINPUT89), .Z(n821) );
  NAND2_X1 U876 ( .A1(n876), .A2(G104), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G140), .A2(n610), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n786), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G128), .A2(n879), .ZN(n788) );
  NAND2_X1 U881 ( .A1(G116), .A2(n880), .ZN(n787) );
  NAND2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U883 ( .A(KEYINPUT90), .B(n789), .Z(n790) );
  XNOR2_X1 U884 ( .A(KEYINPUT35), .B(n790), .ZN(n791) );
  NOR2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n793), .ZN(n896) );
  OR2_X1 U887 ( .A1(n821), .A2(n896), .ZN(n819) );
  NAND2_X1 U888 ( .A1(n794), .A2(n819), .ZN(n920) );
  NAND2_X1 U889 ( .A1(n823), .A2(n920), .ZN(n808) );
  AND2_X1 U890 ( .A1(n989), .A2(n808), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n975), .A2(KEYINPUT33), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n518), .A2(n520), .ZN(n810) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n797) );
  XOR2_X1 U894 ( .A(n797), .B(KEYINPUT24), .Z(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U896 ( .A(KEYINPUT95), .B(n800), .Z(n807) );
  NAND2_X1 U897 ( .A1(G166), .A2(G8), .ZN(n801) );
  NOR2_X1 U898 ( .A1(G2090), .A2(n801), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n808), .A2(n514), .ZN(n809) );
  XNOR2_X1 U902 ( .A(n811), .B(KEYINPUT105), .ZN(n813) );
  XNOR2_X1 U903 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U904 ( .A1(n971), .A2(n823), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n826) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n891), .ZN(n928) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n887), .ZN(n921) );
  NOR2_X1 U909 ( .A1(n814), .A2(n921), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U911 ( .A1(n928), .A2(n817), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n821), .A2(n896), .ZN(n940) );
  NAND2_X1 U915 ( .A1(n822), .A2(n940), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U918 ( .A(n828), .B(n827), .ZN(G329) );
  NAND2_X1 U919 ( .A1(n829), .A2(G2106), .ZN(n830) );
  XOR2_X1 U920 ( .A(KEYINPUT107), .B(n830), .Z(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U931 ( .A(G1956), .B(KEYINPUT41), .ZN(n845) );
  XOR2_X1 U932 ( .A(G1971), .B(G1961), .Z(n837) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1976), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(G1966), .B(G1981), .Z(n839) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT108), .B(G2474), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(G227) );
  NAND2_X1 U951 ( .A1(n876), .A2(G100), .ZN(n854) );
  XOR2_X1 U952 ( .A(KEYINPUT109), .B(n854), .Z(n856) );
  NAND2_X1 U953 ( .A1(n880), .A2(G112), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT110), .B(n857), .ZN(n862) );
  NAND2_X1 U956 ( .A1(G124), .A2(n879), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G136), .A2(n610), .ZN(n859) );
  NAND2_X1 U959 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(G162) );
  XNOR2_X1 U961 ( .A(n925), .B(G162), .ZN(n895) );
  NAND2_X1 U962 ( .A1(n876), .A2(G106), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n863), .B(KEYINPUT112), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G142), .A2(n610), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT45), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G118), .A2(n880), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G130), .A2(n879), .ZN(n869) );
  XNOR2_X1 U970 ( .A(KEYINPUT111), .B(n869), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n875) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT115), .B(KEYINPUT113), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n889) );
  NAND2_X1 U976 ( .A1(n876), .A2(G103), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G139), .A2(n610), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n886) );
  NAND2_X1 U979 ( .A1(G127), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G115), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n883), .Z(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT47), .B(n884), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n933) );
  XNOR2_X1 U985 ( .A(n887), .B(n933), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(G160), .B(n890), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n891), .B(G164), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n969), .B(G286), .ZN(n900) );
  XNOR2_X1 U994 ( .A(G171), .B(n981), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  XNOR2_X1 U998 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n916) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2430), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G2438), .B(G2443), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n913) );
  XOR2_X1 U1004 ( .A(G2435), .B(G2454), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G1341), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1007 ( .A(G2446), .B(G2427), .Z(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n914), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n919), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G171), .ZN(G301) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(G160), .B(G2084), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT117), .B(n926), .ZN(n931) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT51), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT118), .B(n932), .Z(n938) );
  XOR2_X1 U1029 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n936), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n941), .B(KEYINPUT119), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n942), .ZN(n943) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n964), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1040 ( .A(G34), .B(KEYINPUT121), .Z(n946) );
  XNOR2_X1 U1041 ( .A(G2084), .B(KEYINPUT54), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(n946), .B(n945), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n962) );
  XOR2_X1 U1045 ( .A(G2067), .B(G26), .Z(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G2072), .B(G33), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n952), .B(G27), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(n959), .B(KEYINPUT120), .Z(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n966) );
  INV_X1 U1059 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n967), .ZN(n1024) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1063 ( .A(n968), .B(G1956), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G1341), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n987) );
  XNOR2_X1 U1067 ( .A(G166), .B(G1971), .ZN(n974) );
  XOR2_X1 U1068 ( .A(KEYINPUT124), .B(n974), .Z(n977) );
  XOR2_X1 U1069 ( .A(n975), .B(KEYINPUT123), .Z(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT125), .ZN(n985) );
  XOR2_X1 U1073 ( .A(G1348), .B(n981), .Z(n983) );
  XOR2_X1 U1074 ( .A(G171), .B(G1961), .Z(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(KEYINPUT126), .B(n988), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(KEYINPUT57), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n992), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1022) );
  INV_X1 U1085 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1086 ( .A(KEYINPUT127), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(G5), .ZN(n1010) );
  XNOR2_X1 U1088 ( .A(G20), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(G1976), .B(G23), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

