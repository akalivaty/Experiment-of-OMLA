//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G134gat), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n207), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n207), .B2(new_n215), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT2), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(new_n235), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n217), .A2(new_n218), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n225), .A2(new_n235), .ZN(new_n238));
  INV_X1    g037(.A(new_n216), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT66), .B1(new_n212), .B2(new_n214), .ZN(new_n240));
  AOI211_X1 g039(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n209), .C2(new_n211), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n207), .A2(new_n215), .A3(new_n216), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n204), .B1(new_n237), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT77), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n247), .B(new_n204), .C1(new_n237), .C2(new_n244), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(KEYINPUT5), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n246), .A2(KEYINPUT78), .A3(KEYINPUT5), .A4(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n225), .A2(new_n235), .A3(KEYINPUT75), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n254), .A2(new_n242), .A3(new_n243), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n243), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n203), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n252), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n260), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n275), .A4(new_n203), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n271), .A2(new_n272), .A3(new_n275), .A4(new_n268), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n204), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G57gat), .B(G85gat), .Z(new_n282));
  XNOR2_X1  g081(.A(G1gat), .B(G29gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n281), .A2(KEYINPUT6), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n290), .B(new_n286), .C1(new_n270), .C2(new_n280), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n286), .A3(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT81), .B1(new_n281), .B2(new_n287), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n289), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT64), .B1(new_n308), .B2(KEYINPUT23), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n308), .B2(KEYINPUT23), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n307), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT27), .B(G183gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n304), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n314), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n330), .A3(new_n304), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n325), .A2(new_n329), .A3(new_n299), .A4(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n301), .A2(new_n305), .A3(new_n318), .A4(new_n302), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n333), .A2(new_n314), .A3(new_n334), .A4(new_n309), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT25), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n322), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G226gat), .ZN(new_n339));
  INV_X1    g138(.A(G233gat), .ZN(new_n340));
  OAI22_X1  g139(.A1(new_n338), .A2(KEYINPUT29), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n332), .A2(new_n336), .ZN(new_n342));
  NOR4_X1   g141(.A1(new_n311), .A2(new_n315), .A3(new_n312), .A4(KEYINPUT25), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n306), .B1(new_n343), .B2(new_n320), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(G226gat), .A3(G233gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(G197gat), .A2(G204gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT22), .ZN(new_n350));
  NAND2_X1  g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n355));
  NOR2_X1   g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n352), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n349), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n351), .A2(new_n350), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n355), .A3(new_n351), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT73), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n341), .B(new_n346), .C1(new_n366), .C2(new_n367), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n374), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n374), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n380), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n202), .B1(new_n298), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n281), .A2(KEYINPUT81), .A3(new_n287), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n293), .A3(new_n292), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n288), .B1(new_n387), .B2(new_n296), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n389));
  XNOR2_X1  g188(.A(G22gat), .B(G50gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n266), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n368), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n254), .A2(new_n255), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n359), .B2(new_n365), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n392), .B1(new_n366), .B2(new_n367), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT83), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n392), .C1(new_n366), .C2(new_n367), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n265), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n236), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT84), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n407), .A3(new_n236), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n394), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n395), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n399), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT31), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  AOI211_X1 g214(.A(new_n413), .B(new_n399), .C1(new_n409), .C2(new_n410), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n391), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT3), .B1(new_n400), .B2(KEYINPUT83), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT84), .B(new_n238), .C1(new_n418), .C2(new_n403), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n407), .B1(new_n404), .B2(new_n236), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n395), .B1(new_n421), .B2(new_n394), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n413), .B1(new_n422), .B2(new_n399), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n411), .A2(new_n414), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n390), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n417), .A2(KEYINPUT85), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n415), .A2(new_n416), .A3(new_n391), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n390), .B1(new_n423), .B2(new_n424), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n385), .A2(new_n389), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n281), .A2(KEYINPUT87), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n270), .A2(new_n433), .A3(new_n280), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n287), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n294), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n289), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n380), .A2(KEYINPUT37), .A3(new_n381), .ZN(new_n438));
  INV_X1    g237(.A(new_n378), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n440));
  AOI21_X1  g239(.A(new_n373), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n442), .A2(KEYINPUT38), .B1(new_n373), .B2(new_n439), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT38), .B1(new_n378), .B2(KEYINPUT37), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n273), .A2(new_n204), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n237), .A2(new_n244), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(KEYINPUT39), .C1(new_n204), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n450), .A2(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(KEYINPUT86), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n273), .A2(new_n204), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n449), .A2(KEYINPUT40), .A3(new_n286), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT88), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n286), .A3(new_n453), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT40), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n384), .A2(new_n455), .A3(new_n435), .A4(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n428), .A2(new_n429), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n446), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n217), .A2(new_n218), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n342), .A2(new_n464), .A3(new_n344), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n264), .B1(new_n322), .B2(new_n337), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT32), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n467), .B2(KEYINPUT33), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n467), .A2(new_n471), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT69), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT69), .ZN(new_n484));
  NOR4_X1   g283(.A1(new_n467), .A2(new_n484), .A3(new_n471), .A4(new_n481), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n473), .A2(new_n478), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n466), .A3(new_n463), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT34), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n478), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n472), .A3(new_n469), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n488), .C1(new_n483), .C2(new_n485), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(KEYINPUT70), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n486), .A2(new_n495), .A3(new_n489), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n462), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n490), .A2(new_n493), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(new_n462), .ZN(new_n500));
  AOI211_X1 g299(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n490), .C2(new_n493), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n431), .A2(new_n461), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n417), .A2(new_n425), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n383), .A2(new_n490), .A3(new_n493), .ZN(new_n505));
  NOR4_X1   g304(.A1(new_n504), .A2(new_n505), .A3(new_n437), .A4(KEYINPUT35), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n494), .A2(new_n496), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n507), .A2(new_n425), .A3(new_n417), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n385), .A2(new_n508), .A3(new_n389), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT90), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n512));
  INV_X1    g311(.A(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n430), .A2(new_n426), .ZN(new_n515));
  INV_X1    g314(.A(new_n389), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT82), .B1(new_n388), .B2(new_n383), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n446), .A2(new_n459), .A3(new_n460), .ZN(new_n519));
  INV_X1    g318(.A(new_n502), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(G29gat), .A2(G36gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G43gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G50gat), .ZN(new_n532));
  INV_X1    g331(.A(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G43gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT15), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n534), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT92), .B(G50gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(new_n531), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT93), .B1(new_n539), .B2(KEYINPUT15), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(KEYINPUT92), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G50gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n543), .A3(new_n531), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n534), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n528), .A2(KEYINPUT94), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n529), .B1(new_n535), .B2(KEYINPUT91), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n532), .A2(new_n534), .A3(new_n552), .A4(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n526), .A2(new_n527), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n550), .A2(new_n551), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n536), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT95), .B(KEYINPUT17), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n561), .A2(G1gat), .ZN(new_n562));
  INV_X1    g361(.A(G8gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n561), .B1(new_n564), .B2(G1gat), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n562), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n536), .B(KEYINPUT17), .C1(new_n549), .C2(new_n557), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n560), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n558), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n571), .B(new_n558), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n573), .B(KEYINPUT13), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n570), .A2(KEYINPUT18), .A3(new_n572), .A4(new_n573), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  INV_X1    g381(.A(G197gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT11), .B(G169gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT12), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n581), .A2(KEYINPUT96), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT96), .B1(new_n581), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n576), .A2(new_n579), .A3(new_n580), .A4(new_n587), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT98), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n581), .A2(new_n588), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n581), .A2(KEYINPUT96), .A3(new_n588), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n592), .B(KEYINPUT97), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT101), .B(G85gat), .ZN(new_n606));
  INV_X1    g405(.A(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT7), .ZN(new_n610));
  INV_X1    g409(.A(G99gat), .ZN(new_n611));
  INV_X1    g410(.A(G106gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT8), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G99gat), .B(G106gat), .Z(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n560), .B(new_n569), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n616), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n558), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n625), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G57gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G64gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(G71gat), .A2(G78gat), .ZN(new_n634));
  OR2_X1    g433(.A1(G71gat), .A2(G78gat), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT9), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n635), .A2(new_n634), .ZN(new_n638));
  OR2_X1    g437(.A1(G57gat), .A2(G64gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(G57gat), .A2(G64gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(KEYINPUT9), .A3(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n633), .A2(new_n637), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n568), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G183gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n568), .A2(new_n303), .A3(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G211gat), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  XNOR2_X1  g455(.A(G127gat), .B(G155gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n653), .B2(new_n654), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G230gat), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n340), .ZN(new_n663));
  INV_X1    g462(.A(new_n642), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n617), .B2(new_n616), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n614), .A2(new_n615), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n614), .A2(new_n615), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n642), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n619), .A2(KEYINPUT10), .A3(new_n642), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n663), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n665), .A2(new_n668), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(G176gat), .B(G204gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n673), .A2(new_n675), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n630), .A2(new_n661), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT103), .Z(new_n685));
  NAND4_X1  g484(.A1(new_n511), .A2(new_n523), .A3(new_n605), .A4(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n298), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g488(.A1(new_n686), .A2(new_n383), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n564), .A2(new_n563), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n690), .A2(new_n691), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G8gat), .B1(new_n686), .B2(new_n383), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n686), .A2(new_n383), .A3(new_n692), .A4(new_n694), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n696), .B(new_n702), .C1(new_n698), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1325gat));
  INV_X1    g503(.A(G15gat), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n686), .A2(new_n705), .A3(new_n520), .ZN(new_n706));
  INV_X1    g505(.A(new_n499), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n705), .B2(new_n708), .ZN(G1326gat));
  INV_X1    g508(.A(new_n515), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n686), .A2(G22gat), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G22gat), .B1(new_n686), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n630), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n511), .A2(new_n523), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n385), .A2(new_n389), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n502), .B1(new_n719), .B2(new_n515), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n519), .A2(new_n720), .B1(new_n512), .B2(new_n513), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n716), .B1(new_n721), .B2(new_n630), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n600), .A2(new_n601), .ZN(new_n723));
  INV_X1    g522(.A(new_n683), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n661), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT106), .Z(new_n727));
  NAND3_X1  g526(.A1(new_n718), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n388), .ZN(new_n729));
  AND4_X1   g528(.A1(new_n511), .A2(new_n523), .A3(new_n605), .A4(new_n725), .ZN(new_n730));
  INV_X1    g529(.A(G29gat), .ZN(new_n731));
  INV_X1    g530(.A(new_n630), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n298), .A4(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(KEYINPUT45), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(KEYINPUT45), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n729), .B1(new_n734), .B2(new_n735), .ZN(G1328gat));
  AND2_X1   g535(.A1(new_n730), .A2(new_n732), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n383), .A2(G36gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  OAI21_X1  g539(.A(G36gat), .B1(new_n728), .B2(new_n383), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n737), .A2(new_n742), .A3(new_n738), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(G1329gat));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n722), .A3(new_n502), .A4(new_n727), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G43gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n531), .A3(new_n707), .A4(new_n732), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT47), .B1(new_n748), .B2(KEYINPUT107), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n750), .B(new_n751), .C1(new_n746), .C2(new_n747), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n752), .ZN(G1330gat));
  OAI21_X1  g552(.A(new_n538), .B1(new_n728), .B2(new_n460), .ZN(new_n754));
  INV_X1    g553(.A(new_n538), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n730), .A2(new_n515), .A3(new_n755), .A4(new_n732), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT48), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n538), .B1(new_n728), .B2(new_n710), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT108), .A4(KEYINPUT48), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n514), .A2(new_n521), .ZN(new_n766));
  INV_X1    g565(.A(new_n661), .ZN(new_n767));
  NOR4_X1   g566(.A1(new_n723), .A2(new_n732), .A3(new_n767), .A4(new_n683), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT109), .Z(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n388), .B(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g573(.A(new_n383), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n777), .B(new_n778), .Z(G1333gat));
  NAND3_X1  g578(.A1(new_n771), .A2(G71gat), .A3(new_n502), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n770), .A2(new_n499), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(G71gat), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n771), .A2(new_n515), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n723), .A2(new_n661), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n718), .A2(new_n722), .A3(new_n724), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n388), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n766), .A2(new_n732), .A3(new_n787), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n766), .A2(KEYINPUT51), .A3(new_n732), .A4(new_n787), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n724), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n298), .A2(new_n606), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n789), .A2(new_n606), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n788), .B2(new_n383), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n384), .A2(new_n607), .A3(new_n724), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n804), .A3(KEYINPUT52), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n798), .B(new_n803), .C1(new_n799), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n788), .B2(new_n520), .ZN(new_n809));
  INV_X1    g608(.A(new_n794), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n499), .A2(G99gat), .A3(new_n683), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT115), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(G1338gat));
  OAI21_X1  g612(.A(G106gat), .B1(new_n788), .B2(new_n460), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n794), .A2(new_n612), .A3(new_n504), .A4(new_n724), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G106gat), .B1(new_n788), .B2(new_n710), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n815), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(new_n816), .ZN(G1339gat));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n672), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n822), .B2(new_n679), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n824), .B(new_n681), .C1(new_n672), .C2(new_n821), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n670), .A2(new_n671), .A3(new_n663), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n673), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT55), .B(new_n828), .C1(new_n823), .C2(new_n825), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n682), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(KEYINPUT117), .A3(new_n682), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n577), .A2(new_n578), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n573), .B1(new_n570), .B2(new_n572), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n586), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n601), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n835), .B(new_n732), .C1(KEYINPUT118), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n601), .B2(new_n838), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n601), .A2(new_n838), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n835), .A2(new_n723), .B1(new_n843), .B2(new_n724), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n840), .A2(new_n842), .B1(new_n844), .B2(new_n732), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n767), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n684), .A2(new_n723), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n849), .A2(new_n383), .A3(new_n772), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n508), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n210), .A3(new_n723), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n847), .B1(new_n845), .B2(new_n767), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n515), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n854), .A2(new_n298), .A3(new_n383), .A4(new_n707), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n604), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n851), .A2(new_n208), .A3(new_n724), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n855), .B2(new_n683), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n855), .A2(new_n861), .A3(new_n767), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n851), .A2(new_n661), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT119), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n861), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n866), .A3(new_n732), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n855), .B2(new_n630), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n502), .A2(new_n460), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n850), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(new_n226), .A3(new_n605), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n853), .A2(KEYINPUT57), .A3(new_n460), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n829), .A2(new_n831), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n595), .A2(new_n603), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n843), .A2(new_n724), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n732), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n732), .B1(new_n839), .B2(KEYINPUT118), .ZN(new_n880));
  INV_X1    g679(.A(new_n829), .ZN(new_n881));
  INV_X1    g680(.A(new_n834), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT117), .B1(new_n830), .B2(new_n682), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n880), .A2(new_n884), .A3(new_n842), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n767), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n848), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n710), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n502), .A2(new_n388), .A3(new_n384), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n875), .A2(new_n888), .A3(new_n723), .A4(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n874), .B1(G141gat), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n888), .A3(new_n889), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n604), .ZN(new_n894));
  XNOR2_X1  g693(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n891), .A2(new_n892), .B1(new_n896), .B2(new_n874), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n873), .A2(new_n228), .A3(new_n724), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n685), .A2(new_n604), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n886), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n710), .A2(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n900), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT57), .B1(new_n853), .B2(new_n460), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n724), .A3(new_n889), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n899), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n899), .B(G148gat), .C1(new_n893), .C2(new_n683), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n898), .B1(new_n911), .B2(new_n913), .ZN(G1345gat));
  AOI21_X1  g713(.A(G155gat), .B1(new_n873), .B2(new_n661), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n893), .A2(new_n232), .A3(new_n767), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1346gat));
  AOI21_X1  g716(.A(G162gat), .B1(new_n873), .B2(new_n732), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n893), .A2(new_n233), .A3(new_n630), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1347gat));
  AND4_X1   g719(.A1(new_n388), .A2(new_n849), .A3(new_n384), .A4(new_n508), .ZN(new_n921));
  INV_X1    g720(.A(G169gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n723), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n772), .A2(new_n383), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n854), .A2(new_n707), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n605), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT122), .B1(new_n927), .B2(G169gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  AOI21_X1  g729(.A(G176gat), .B1(new_n921), .B2(new_n724), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n925), .A2(new_n683), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(G176gat), .B2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n925), .B2(new_n767), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n921), .A2(new_n323), .A3(new_n661), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n936), .B(new_n937), .Z(G1350gat));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n304), .A3(new_n732), .ZN(new_n939));
  OAI21_X1  g738(.A(G190gat), .B1(new_n925), .B2(new_n630), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n520), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n908), .A2(new_n604), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(G197gat), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n872), .ZN(new_n949));
  NOR4_X1   g748(.A1(new_n853), .A2(new_n298), .A3(new_n949), .A4(new_n383), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n583), .A3(new_n723), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT124), .Z(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n954), .A3(new_n724), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g755(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n908), .A2(new_n683), .A3(new_n944), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n954), .B2(new_n959), .ZN(G1353gat));
  INV_X1    g759(.A(G211gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n950), .A2(new_n961), .A3(new_n661), .ZN(new_n962));
  INV_X1    g761(.A(new_n944), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n906), .A2(new_n661), .A3(new_n907), .A4(new_n963), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n962), .B(new_n969), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1354gat));
  AND4_X1   g770(.A1(G218gat), .A2(new_n909), .A3(new_n732), .A4(new_n963), .ZN(new_n972));
  AOI21_X1  g771(.A(G218gat), .B1(new_n950), .B2(new_n732), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


